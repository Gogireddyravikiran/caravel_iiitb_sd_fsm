magic
tech sky130B
magscale 1 2
timestamp 1662965032
<< obsli1 >>
rect 1104 2159 8832 7633
<< obsm1 >>
rect 14 2128 9738 7664
<< metal2 >>
rect 18 9200 74 10000
rect 9678 9200 9734 10000
rect 18 0 74 800
rect 9678 0 9734 800
<< obsm2 >>
rect 130 9144 9622 9200
rect 20 856 9732 9144
rect 130 800 9622 856
<< obsm3 >>
rect 1920 2143 8080 7649
<< metal4 >>
rect 1918 2128 2238 7664
rect 2892 2128 3212 7664
rect 3866 2128 4186 7664
rect 4840 2128 5160 7664
rect 5814 2128 6134 7664
rect 6788 2128 7108 7664
rect 7762 2128 8082 7664
<< labels >>
rlabel metal2 s 18 0 74 800 6 clock
port 1 nsew signal input
rlabel metal2 s 18 9200 74 10000 6 detector_out
port 2 nsew signal output
rlabel metal2 s 9678 9200 9734 10000 6 reset
port 3 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 sequence_in
port 4 nsew signal input
rlabel metal4 s 1918 2128 2238 7664 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 3866 2128 4186 7664 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 5814 2128 6134 7664 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 7762 2128 8082 7664 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 2892 2128 3212 7664 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 4840 2128 5160 7664 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 6788 2128 7108 7664 6 vssd1
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 192282
string GDS_FILE /home/ravi/Desktop/caravel_iiitb_sd_fsm/openlane/iiitb_sd_fsm/runs/22_09_12_12_12/results/signoff/iiitb_sd_fsm.magic.gds
string GDS_START 106888
<< end >>

