magic
tech sky130B
magscale 1 2
timestamp 1662965030
<< viali >>
rect 1501 7497 1535 7531
rect 1685 7361 1719 7395
rect 7849 7293 7883 7327
rect 8125 7293 8159 7327
rect 8125 6817 8159 6851
rect 4353 5661 4387 5695
rect 6745 5661 6779 5695
rect 4629 5593 4663 5627
rect 6653 5593 6687 5627
rect 6101 5525 6135 5559
rect 4261 5321 4295 5355
rect 3893 5253 3927 5287
rect 2789 5185 2823 5219
rect 3709 5185 3743 5219
rect 3985 5185 4019 5219
rect 4077 5185 4111 5219
rect 4905 5185 4939 5219
rect 7481 5185 7515 5219
rect 3249 5117 3283 5151
rect 2881 4981 2915 5015
rect 4721 4981 4755 5015
rect 7389 4981 7423 5015
rect 3065 4777 3099 4811
rect 3801 4777 3835 4811
rect 4169 4777 4203 4811
rect 4905 4777 4939 4811
rect 3249 4709 3283 4743
rect 4813 4641 4847 4675
rect 7941 4641 7975 4675
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 4997 4573 5031 4607
rect 5089 4573 5123 4607
rect 5549 4573 5583 4607
rect 6193 4573 6227 4607
rect 2881 4505 2915 4539
rect 6469 4505 6503 4539
rect 3091 4437 3125 4471
rect 5733 4437 5767 4471
rect 3433 4233 3467 4267
rect 6377 4233 6411 4267
rect 6561 4165 6595 4199
rect 3525 4097 3559 4131
rect 4169 4097 4203 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5825 4097 5859 4131
rect 6929 3961 6963 3995
rect 3985 3893 4019 3927
rect 5733 3893 5767 3927
rect 6561 3893 6595 3927
rect 6101 3689 6135 3723
rect 4353 3485 4387 3519
rect 4629 3417 4663 3451
rect 3801 3009 3835 3043
rect 3709 2941 3743 2975
rect 4169 2941 4203 2975
rect 1593 2601 1627 2635
rect 7941 2601 7975 2635
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 7481 2397 7515 2431
rect 8125 2397 8159 2431
<< metal1 >>
rect 1104 7642 8832 7664
rect 1104 7590 2898 7642
rect 2950 7590 2962 7642
rect 3014 7590 3026 7642
rect 3078 7590 3090 7642
rect 3142 7590 3154 7642
rect 3206 7590 4846 7642
rect 4898 7590 4910 7642
rect 4962 7590 4974 7642
rect 5026 7590 5038 7642
rect 5090 7590 5102 7642
rect 5154 7590 6794 7642
rect 6846 7590 6858 7642
rect 6910 7590 6922 7642
rect 6974 7590 6986 7642
rect 7038 7590 7050 7642
rect 7102 7590 8832 7642
rect 1104 7568 8832 7590
rect 14 7488 20 7540
rect 72 7528 78 7540
rect 1489 7531 1547 7537
rect 1489 7528 1501 7531
rect 72 7500 1501 7528
rect 72 7488 78 7500
rect 1489 7497 1501 7500
rect 1535 7497 1547 7531
rect 1489 7491 1547 7497
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7524 7296 7849 7324
rect 7524 7284 7530 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 8110 7324 8116 7336
rect 8071 7296 8116 7324
rect 7837 7287 7895 7293
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 1104 7098 8832 7120
rect 1104 7046 1924 7098
rect 1976 7046 1988 7098
rect 2040 7046 2052 7098
rect 2104 7046 2116 7098
rect 2168 7046 2180 7098
rect 2232 7046 3872 7098
rect 3924 7046 3936 7098
rect 3988 7046 4000 7098
rect 4052 7046 4064 7098
rect 4116 7046 4128 7098
rect 4180 7046 5820 7098
rect 5872 7046 5884 7098
rect 5936 7046 5948 7098
rect 6000 7046 6012 7098
rect 6064 7046 6076 7098
rect 6128 7046 7768 7098
rect 7820 7046 7832 7098
rect 7884 7046 7896 7098
rect 7948 7046 7960 7098
rect 8012 7046 8024 7098
rect 8076 7046 8832 7098
rect 1104 7024 8832 7046
rect 8110 6848 8116 6860
rect 8023 6820 8116 6848
rect 8110 6808 8116 6820
rect 8168 6848 8174 6860
rect 9674 6848 9680 6860
rect 8168 6820 9680 6848
rect 8168 6808 8174 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 1104 6554 8832 6576
rect 1104 6502 2898 6554
rect 2950 6502 2962 6554
rect 3014 6502 3026 6554
rect 3078 6502 3090 6554
rect 3142 6502 3154 6554
rect 3206 6502 4846 6554
rect 4898 6502 4910 6554
rect 4962 6502 4974 6554
rect 5026 6502 5038 6554
rect 5090 6502 5102 6554
rect 5154 6502 6794 6554
rect 6846 6502 6858 6554
rect 6910 6502 6922 6554
rect 6974 6502 6986 6554
rect 7038 6502 7050 6554
rect 7102 6502 8832 6554
rect 1104 6480 8832 6502
rect 1104 6010 8832 6032
rect 1104 5958 1924 6010
rect 1976 5958 1988 6010
rect 2040 5958 2052 6010
rect 2104 5958 2116 6010
rect 2168 5958 2180 6010
rect 2232 5958 3872 6010
rect 3924 5958 3936 6010
rect 3988 5958 4000 6010
rect 4052 5958 4064 6010
rect 4116 5958 4128 6010
rect 4180 5958 5820 6010
rect 5872 5958 5884 6010
rect 5936 5958 5948 6010
rect 6000 5958 6012 6010
rect 6064 5958 6076 6010
rect 6128 5958 7768 6010
rect 7820 5958 7832 6010
rect 7884 5958 7896 6010
rect 7948 5958 7960 6010
rect 8012 5958 8024 6010
rect 8076 5958 8832 6010
rect 1104 5936 8832 5958
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 7466 5692 7472 5704
rect 6779 5664 7472 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 4614 5624 4620 5636
rect 4575 5596 4620 5624
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 5842 5596 6653 5624
rect 6641 5593 6653 5596
rect 6687 5593 6699 5627
rect 6641 5587 6699 5593
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6546 5556 6552 5568
rect 6135 5528 6552 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 1104 5466 8832 5488
rect 1104 5414 2898 5466
rect 2950 5414 2962 5466
rect 3014 5414 3026 5466
rect 3078 5414 3090 5466
rect 3142 5414 3154 5466
rect 3206 5414 4846 5466
rect 4898 5414 4910 5466
rect 4962 5414 4974 5466
rect 5026 5414 5038 5466
rect 5090 5414 5102 5466
rect 5154 5414 6794 5466
rect 6846 5414 6858 5466
rect 6910 5414 6922 5466
rect 6974 5414 6986 5466
rect 7038 5414 7050 5466
rect 7102 5414 8832 5466
rect 1104 5392 8832 5414
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4614 5352 4620 5364
rect 4295 5324 4620 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 3881 5287 3939 5293
rect 3881 5253 3893 5287
rect 3927 5284 3939 5287
rect 4706 5284 4712 5296
rect 3927 5256 4712 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 3694 5216 3700 5228
rect 3655 5188 3700 5216
rect 2777 5179 2835 5185
rect 2792 5080 2820 5179
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3844 5188 3985 5216
rect 3844 5176 3850 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 4080 5148 4108 5179
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4304 5188 4905 5216
rect 4304 5176 4310 5188
rect 4893 5185 4905 5188
rect 4939 5185 4951 5219
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 4893 5179 4951 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 3283 5120 4108 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3602 5080 3608 5092
rect 2792 5052 3608 5080
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 1728 4984 2881 5012
rect 1728 4972 1734 4984
rect 2869 4981 2881 4984
rect 2915 5012 2927 5015
rect 4709 5015 4767 5021
rect 4709 5012 4721 5015
rect 2915 4984 4721 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 4709 4981 4721 4984
rect 4755 4981 4767 5015
rect 4709 4975 4767 4981
rect 7377 5015 7435 5021
rect 7377 4981 7389 5015
rect 7423 5012 7435 5015
rect 7466 5012 7472 5024
rect 7423 4984 7472 5012
rect 7423 4981 7435 4984
rect 7377 4975 7435 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 1104 4922 8832 4944
rect 1104 4870 1924 4922
rect 1976 4870 1988 4922
rect 2040 4870 2052 4922
rect 2104 4870 2116 4922
rect 2168 4870 2180 4922
rect 2232 4870 3872 4922
rect 3924 4870 3936 4922
rect 3988 4870 4000 4922
rect 4052 4870 4064 4922
rect 4116 4870 4128 4922
rect 4180 4870 5820 4922
rect 5872 4870 5884 4922
rect 5936 4870 5948 4922
rect 6000 4870 6012 4922
rect 6064 4870 6076 4922
rect 6128 4870 7768 4922
rect 7820 4870 7832 4922
rect 7884 4870 7896 4922
rect 7948 4870 7960 4922
rect 8012 4870 8024 4922
rect 8076 4870 8832 4922
rect 1104 4848 8832 4870
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3510 4808 3516 4820
rect 3099 4780 3516 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 3602 4768 3608 4820
rect 3660 4808 3666 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3660 4780 3801 4808
rect 3660 4768 3666 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 4154 4808 4160 4820
rect 4067 4780 4160 4808
rect 3789 4771 3847 4777
rect 4154 4768 4160 4780
rect 4212 4808 4218 4820
rect 4212 4780 4660 4808
rect 4212 4768 4218 4780
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 4246 4740 4252 4752
rect 3283 4712 4252 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 4632 4740 4660 4780
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4764 4780 4905 4808
rect 4764 4768 4770 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 4632 4712 5120 4740
rect 4614 4672 4620 4684
rect 2884 4644 4620 4672
rect 2884 4545 2912 4644
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4062 4604 4068 4616
rect 3752 4576 4068 4604
rect 3752 4564 3758 4576
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4356 4613 4384 4644
rect 4614 4632 4620 4644
rect 4672 4672 4678 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4672 4644 4813 4672
rect 4672 4632 4678 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 5092 4672 5120 4712
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 5092 4644 7941 4672
rect 5092 4613 5120 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4573 5135 4607
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5077 4567 5135 4573
rect 2869 4539 2927 4545
rect 2869 4505 2881 4539
rect 2915 4505 2927 4539
rect 2869 4499 2927 4505
rect 3786 4496 3792 4548
rect 3844 4536 3850 4548
rect 5000 4536 5028 4567
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 3844 4508 5028 4536
rect 6457 4539 6515 4545
rect 3844 4496 3850 4508
rect 6457 4505 6469 4539
rect 6503 4505 6515 4539
rect 6457 4499 6515 4505
rect 3079 4471 3137 4477
rect 3079 4437 3091 4471
rect 3125 4468 3137 4471
rect 4154 4468 4160 4480
rect 3125 4440 4160 4468
rect 3125 4437 3137 4440
rect 3079 4431 3137 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 5721 4471 5779 4477
rect 5721 4437 5733 4471
rect 5767 4468 5779 4471
rect 6472 4468 6500 4499
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 5767 4440 6500 4468
rect 5767 4437 5779 4440
rect 5721 4431 5779 4437
rect 1104 4378 8832 4400
rect 1104 4326 2898 4378
rect 2950 4326 2962 4378
rect 3014 4326 3026 4378
rect 3078 4326 3090 4378
rect 3142 4326 3154 4378
rect 3206 4326 4846 4378
rect 4898 4326 4910 4378
rect 4962 4326 4974 4378
rect 5026 4326 5038 4378
rect 5090 4326 5102 4378
rect 5154 4326 6794 4378
rect 6846 4326 6858 4378
rect 6910 4326 6922 4378
rect 6974 4326 6986 4378
rect 7038 4326 7050 4378
rect 7102 4326 8832 4378
rect 1104 4304 8832 4326
rect 3421 4267 3479 4273
rect 3421 4233 3433 4267
rect 3467 4264 3479 4267
rect 3786 4264 3792 4276
rect 3467 4236 3792 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 5592 4236 6377 4264
rect 5592 4224 5598 4236
rect 6365 4233 6377 4236
rect 6411 4233 6423 4267
rect 6365 4227 6423 4233
rect 6549 4199 6607 4205
rect 6549 4196 6561 4199
rect 5644 4168 6561 4196
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 4154 4128 4160 4140
rect 4115 4100 4160 4128
rect 3513 4091 3571 4097
rect 3528 4060 3556 4091
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4614 4128 4620 4140
rect 4575 4100 4620 4128
rect 4433 4091 4491 4097
rect 4448 4060 4476 4091
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5644 4060 5672 4168
rect 6549 4165 6561 4168
rect 6595 4196 6607 4199
rect 6638 4196 6644 4208
rect 6595 4168 6644 4196
rect 6595 4165 6607 4168
rect 6549 4159 6607 4165
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 7374 4128 7380 4140
rect 5859 4100 7380 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 3528 4032 5672 4060
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 4062 3992 4068 4004
rect 3844 3964 4068 3992
rect 3844 3952 3850 3964
rect 4062 3952 4068 3964
rect 4120 3992 4126 4004
rect 6914 3992 6920 4004
rect 4120 3964 6592 3992
rect 6875 3964 6920 3992
rect 4120 3952 4126 3964
rect 6564 3936 6592 3964
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3752 3896 3985 3924
rect 3752 3884 3758 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 3973 3887 4031 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 1104 3834 8832 3856
rect 1104 3782 1924 3834
rect 1976 3782 1988 3834
rect 2040 3782 2052 3834
rect 2104 3782 2116 3834
rect 2168 3782 2180 3834
rect 2232 3782 3872 3834
rect 3924 3782 3936 3834
rect 3988 3782 4000 3834
rect 4052 3782 4064 3834
rect 4116 3782 4128 3834
rect 4180 3782 5820 3834
rect 5872 3782 5884 3834
rect 5936 3782 5948 3834
rect 6000 3782 6012 3834
rect 6064 3782 6076 3834
rect 6128 3782 7768 3834
rect 7820 3782 7832 3834
rect 7884 3782 7896 3834
rect 7948 3782 7960 3834
rect 8012 3782 8024 3834
rect 8076 3782 8832 3834
rect 1104 3760 8832 3782
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 4672 3692 6101 3720
rect 4672 3680 4678 3692
rect 6089 3689 6101 3692
rect 6135 3720 6147 3723
rect 6914 3720 6920 3732
rect 6135 3692 6920 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 6178 3584 6184 3596
rect 4356 3556 6184 3584
rect 4356 3528 4384 3556
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 4338 3516 4344 3528
rect 4299 3488 4344 3516
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 4212 3420 4629 3448
rect 4212 3408 4218 3420
rect 4617 3417 4629 3420
rect 4663 3417 4675 3451
rect 4617 3411 4675 3417
rect 1104 3290 8832 3312
rect 1104 3238 2898 3290
rect 2950 3238 2962 3290
rect 3014 3238 3026 3290
rect 3078 3238 3090 3290
rect 3142 3238 3154 3290
rect 3206 3238 4846 3290
rect 4898 3238 4910 3290
rect 4962 3238 4974 3290
rect 5026 3238 5038 3290
rect 5090 3238 5102 3290
rect 5154 3238 6794 3290
rect 6846 3238 6858 3290
rect 6910 3238 6922 3290
rect 6974 3238 6986 3290
rect 7038 3238 7050 3290
rect 7102 3238 8832 3290
rect 1104 3216 8832 3238
rect 3786 3040 3792 3052
rect 3747 3012 3792 3040
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 3694 2972 3700 2984
rect 3655 2944 3700 2972
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 4154 2972 4160 2984
rect 4115 2944 4160 2972
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 9674 2836 9680 2848
rect 8168 2808 9680 2836
rect 8168 2796 8174 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 1104 2746 8832 2768
rect 1104 2694 1924 2746
rect 1976 2694 1988 2746
rect 2040 2694 2052 2746
rect 2104 2694 2116 2746
rect 2168 2694 2180 2746
rect 2232 2694 3872 2746
rect 3924 2694 3936 2746
rect 3988 2694 4000 2746
rect 4052 2694 4064 2746
rect 4116 2694 4128 2746
rect 4180 2694 5820 2746
rect 5872 2694 5884 2746
rect 5936 2694 5948 2746
rect 6000 2694 6012 2746
rect 6064 2694 6076 2746
rect 6128 2694 7768 2746
rect 7820 2694 7832 2746
rect 7884 2694 7896 2746
rect 7948 2694 7960 2746
rect 8012 2694 8024 2746
rect 8076 2694 8832 2746
rect 1104 2672 8832 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 4338 2632 4344 2644
rect 1627 2604 4344 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 6972 2604 7941 2632
rect 6972 2592 6978 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2428 1455 2431
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 1443 2400 2053 2428
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 8110 2428 8116 2440
rect 7515 2400 8116 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 1104 2202 8832 2224
rect 1104 2150 2898 2202
rect 2950 2150 2962 2202
rect 3014 2150 3026 2202
rect 3078 2150 3090 2202
rect 3142 2150 3154 2202
rect 3206 2150 4846 2202
rect 4898 2150 4910 2202
rect 4962 2150 4974 2202
rect 5026 2150 5038 2202
rect 5090 2150 5102 2202
rect 5154 2150 6794 2202
rect 6846 2150 6858 2202
rect 6910 2150 6922 2202
rect 6974 2150 6986 2202
rect 7038 2150 7050 2202
rect 7102 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 2898 7590 2950 7642
rect 2962 7590 3014 7642
rect 3026 7590 3078 7642
rect 3090 7590 3142 7642
rect 3154 7590 3206 7642
rect 4846 7590 4898 7642
rect 4910 7590 4962 7642
rect 4974 7590 5026 7642
rect 5038 7590 5090 7642
rect 5102 7590 5154 7642
rect 6794 7590 6846 7642
rect 6858 7590 6910 7642
rect 6922 7590 6974 7642
rect 6986 7590 7038 7642
rect 7050 7590 7102 7642
rect 20 7488 72 7540
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 7472 7284 7524 7336
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 1924 7046 1976 7098
rect 1988 7046 2040 7098
rect 2052 7046 2104 7098
rect 2116 7046 2168 7098
rect 2180 7046 2232 7098
rect 3872 7046 3924 7098
rect 3936 7046 3988 7098
rect 4000 7046 4052 7098
rect 4064 7046 4116 7098
rect 4128 7046 4180 7098
rect 5820 7046 5872 7098
rect 5884 7046 5936 7098
rect 5948 7046 6000 7098
rect 6012 7046 6064 7098
rect 6076 7046 6128 7098
rect 7768 7046 7820 7098
rect 7832 7046 7884 7098
rect 7896 7046 7948 7098
rect 7960 7046 8012 7098
rect 8024 7046 8076 7098
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 9680 6808 9732 6860
rect 2898 6502 2950 6554
rect 2962 6502 3014 6554
rect 3026 6502 3078 6554
rect 3090 6502 3142 6554
rect 3154 6502 3206 6554
rect 4846 6502 4898 6554
rect 4910 6502 4962 6554
rect 4974 6502 5026 6554
rect 5038 6502 5090 6554
rect 5102 6502 5154 6554
rect 6794 6502 6846 6554
rect 6858 6502 6910 6554
rect 6922 6502 6974 6554
rect 6986 6502 7038 6554
rect 7050 6502 7102 6554
rect 1924 5958 1976 6010
rect 1988 5958 2040 6010
rect 2052 5958 2104 6010
rect 2116 5958 2168 6010
rect 2180 5958 2232 6010
rect 3872 5958 3924 6010
rect 3936 5958 3988 6010
rect 4000 5958 4052 6010
rect 4064 5958 4116 6010
rect 4128 5958 4180 6010
rect 5820 5958 5872 6010
rect 5884 5958 5936 6010
rect 5948 5958 6000 6010
rect 6012 5958 6064 6010
rect 6076 5958 6128 6010
rect 7768 5958 7820 6010
rect 7832 5958 7884 6010
rect 7896 5958 7948 6010
rect 7960 5958 8012 6010
rect 8024 5958 8076 6010
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 7472 5652 7524 5704
rect 4620 5627 4672 5636
rect 4620 5593 4629 5627
rect 4629 5593 4663 5627
rect 4663 5593 4672 5627
rect 4620 5584 4672 5593
rect 6552 5516 6604 5568
rect 2898 5414 2950 5466
rect 2962 5414 3014 5466
rect 3026 5414 3078 5466
rect 3090 5414 3142 5466
rect 3154 5414 3206 5466
rect 4846 5414 4898 5466
rect 4910 5414 4962 5466
rect 4974 5414 5026 5466
rect 5038 5414 5090 5466
rect 5102 5414 5154 5466
rect 6794 5414 6846 5466
rect 6858 5414 6910 5466
rect 6922 5414 6974 5466
rect 6986 5414 7038 5466
rect 7050 5414 7102 5466
rect 4620 5312 4672 5364
rect 4712 5244 4764 5296
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3792 5176 3844 5228
rect 4252 5176 4304 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 3608 5040 3660 5092
rect 1676 4972 1728 5024
rect 7472 4972 7524 5024
rect 1924 4870 1976 4922
rect 1988 4870 2040 4922
rect 2052 4870 2104 4922
rect 2116 4870 2168 4922
rect 2180 4870 2232 4922
rect 3872 4870 3924 4922
rect 3936 4870 3988 4922
rect 4000 4870 4052 4922
rect 4064 4870 4116 4922
rect 4128 4870 4180 4922
rect 5820 4870 5872 4922
rect 5884 4870 5936 4922
rect 5948 4870 6000 4922
rect 6012 4870 6064 4922
rect 6076 4870 6128 4922
rect 7768 4870 7820 4922
rect 7832 4870 7884 4922
rect 7896 4870 7948 4922
rect 7960 4870 8012 4922
rect 8024 4870 8076 4922
rect 3516 4768 3568 4820
rect 3608 4768 3660 4820
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 4252 4700 4304 4752
rect 4712 4768 4764 4820
rect 3700 4564 3752 4616
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 4620 4632 4672 4684
rect 5540 4607 5592 4616
rect 3792 4496 3844 4548
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 4160 4428 4212 4480
rect 7472 4496 7524 4548
rect 2898 4326 2950 4378
rect 2962 4326 3014 4378
rect 3026 4326 3078 4378
rect 3090 4326 3142 4378
rect 3154 4326 3206 4378
rect 4846 4326 4898 4378
rect 4910 4326 4962 4378
rect 4974 4326 5026 4378
rect 5038 4326 5090 4378
rect 5102 4326 5154 4378
rect 6794 4326 6846 4378
rect 6858 4326 6910 4378
rect 6922 4326 6974 4378
rect 6986 4326 7038 4378
rect 7050 4326 7102 4378
rect 3792 4224 3844 4276
rect 5540 4224 5592 4276
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 6644 4156 6696 4208
rect 7380 4088 7432 4140
rect 3792 3952 3844 4004
rect 4068 3952 4120 4004
rect 6920 3995 6972 4004
rect 6920 3961 6929 3995
rect 6929 3961 6963 3995
rect 6963 3961 6972 3995
rect 6920 3952 6972 3961
rect 3700 3884 3752 3936
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 1924 3782 1976 3834
rect 1988 3782 2040 3834
rect 2052 3782 2104 3834
rect 2116 3782 2168 3834
rect 2180 3782 2232 3834
rect 3872 3782 3924 3834
rect 3936 3782 3988 3834
rect 4000 3782 4052 3834
rect 4064 3782 4116 3834
rect 4128 3782 4180 3834
rect 5820 3782 5872 3834
rect 5884 3782 5936 3834
rect 5948 3782 6000 3834
rect 6012 3782 6064 3834
rect 6076 3782 6128 3834
rect 7768 3782 7820 3834
rect 7832 3782 7884 3834
rect 7896 3782 7948 3834
rect 7960 3782 8012 3834
rect 8024 3782 8076 3834
rect 4620 3680 4672 3732
rect 6920 3680 6972 3732
rect 6184 3544 6236 3596
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 5724 3476 5776 3528
rect 4160 3408 4212 3460
rect 2898 3238 2950 3290
rect 2962 3238 3014 3290
rect 3026 3238 3078 3290
rect 3090 3238 3142 3290
rect 3154 3238 3206 3290
rect 4846 3238 4898 3290
rect 4910 3238 4962 3290
rect 4974 3238 5026 3290
rect 5038 3238 5090 3290
rect 5102 3238 5154 3290
rect 6794 3238 6846 3290
rect 6858 3238 6910 3290
rect 6922 3238 6974 3290
rect 6986 3238 7038 3290
rect 7050 3238 7102 3290
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 8116 2796 8168 2848
rect 9680 2796 9732 2848
rect 1924 2694 1976 2746
rect 1988 2694 2040 2746
rect 2052 2694 2104 2746
rect 2116 2694 2168 2746
rect 2180 2694 2232 2746
rect 3872 2694 3924 2746
rect 3936 2694 3988 2746
rect 4000 2694 4052 2746
rect 4064 2694 4116 2746
rect 4128 2694 4180 2746
rect 5820 2694 5872 2746
rect 5884 2694 5936 2746
rect 5948 2694 6000 2746
rect 6012 2694 6064 2746
rect 6076 2694 6128 2746
rect 7768 2694 7820 2746
rect 7832 2694 7884 2746
rect 7896 2694 7948 2746
rect 7960 2694 8012 2746
rect 8024 2694 8076 2746
rect 4344 2592 4396 2644
rect 6920 2592 6972 2644
rect 20 2388 72 2440
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 2898 2150 2950 2202
rect 2962 2150 3014 2202
rect 3026 2150 3078 2202
rect 3090 2150 3142 2202
rect 3154 2150 3206 2202
rect 4846 2150 4898 2202
rect 4910 2150 4962 2202
rect 4974 2150 5026 2202
rect 5038 2150 5090 2202
rect 5102 2150 5154 2202
rect 6794 2150 6846 2202
rect 6858 2150 6910 2202
rect 6922 2150 6974 2202
rect 6986 2150 7038 2202
rect 7050 2150 7102 2202
<< metal2 >>
rect 18 9200 74 10000
rect 9678 9200 9734 10000
rect 32 7546 60 9200
rect 2898 7644 3206 7653
rect 2898 7642 2904 7644
rect 2960 7642 2984 7644
rect 3040 7642 3064 7644
rect 3120 7642 3144 7644
rect 3200 7642 3206 7644
rect 2960 7590 2962 7642
rect 3142 7590 3144 7642
rect 2898 7588 2904 7590
rect 2960 7588 2984 7590
rect 3040 7588 3064 7590
rect 3120 7588 3144 7590
rect 3200 7588 3206 7590
rect 2898 7579 3206 7588
rect 4846 7644 5154 7653
rect 4846 7642 4852 7644
rect 4908 7642 4932 7644
rect 4988 7642 5012 7644
rect 5068 7642 5092 7644
rect 5148 7642 5154 7644
rect 4908 7590 4910 7642
rect 5090 7590 5092 7642
rect 4846 7588 4852 7590
rect 4908 7588 4932 7590
rect 4988 7588 5012 7590
rect 5068 7588 5092 7590
rect 5148 7588 5154 7590
rect 4846 7579 5154 7588
rect 6794 7644 7102 7653
rect 6794 7642 6800 7644
rect 6856 7642 6880 7644
rect 6936 7642 6960 7644
rect 7016 7642 7040 7644
rect 7096 7642 7102 7644
rect 6856 7590 6858 7642
rect 7038 7590 7040 7642
rect 6794 7588 6800 7590
rect 6856 7588 6880 7590
rect 6936 7588 6960 7590
rect 7016 7588 7040 7590
rect 7096 7588 7102 7590
rect 6794 7579 7102 7588
rect 20 7540 72 7546
rect 20 7482 72 7488
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1688 5030 1716 7346
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 1924 7100 2232 7109
rect 1924 7098 1930 7100
rect 1986 7098 2010 7100
rect 2066 7098 2090 7100
rect 2146 7098 2170 7100
rect 2226 7098 2232 7100
rect 1986 7046 1988 7098
rect 2168 7046 2170 7098
rect 1924 7044 1930 7046
rect 1986 7044 2010 7046
rect 2066 7044 2090 7046
rect 2146 7044 2170 7046
rect 2226 7044 2232 7046
rect 1924 7035 2232 7044
rect 3872 7100 4180 7109
rect 3872 7098 3878 7100
rect 3934 7098 3958 7100
rect 4014 7098 4038 7100
rect 4094 7098 4118 7100
rect 4174 7098 4180 7100
rect 3934 7046 3936 7098
rect 4116 7046 4118 7098
rect 3872 7044 3878 7046
rect 3934 7044 3958 7046
rect 4014 7044 4038 7046
rect 4094 7044 4118 7046
rect 4174 7044 4180 7046
rect 3872 7035 4180 7044
rect 5820 7100 6128 7109
rect 5820 7098 5826 7100
rect 5882 7098 5906 7100
rect 5962 7098 5986 7100
rect 6042 7098 6066 7100
rect 6122 7098 6128 7100
rect 5882 7046 5884 7098
rect 6064 7046 6066 7098
rect 5820 7044 5826 7046
rect 5882 7044 5906 7046
rect 5962 7044 5986 7046
rect 6042 7044 6066 7046
rect 6122 7044 6128 7046
rect 5820 7035 6128 7044
rect 2898 6556 3206 6565
rect 2898 6554 2904 6556
rect 2960 6554 2984 6556
rect 3040 6554 3064 6556
rect 3120 6554 3144 6556
rect 3200 6554 3206 6556
rect 2960 6502 2962 6554
rect 3142 6502 3144 6554
rect 2898 6500 2904 6502
rect 2960 6500 2984 6502
rect 3040 6500 3064 6502
rect 3120 6500 3144 6502
rect 3200 6500 3206 6502
rect 2898 6491 3206 6500
rect 4846 6556 5154 6565
rect 4846 6554 4852 6556
rect 4908 6554 4932 6556
rect 4988 6554 5012 6556
rect 5068 6554 5092 6556
rect 5148 6554 5154 6556
rect 4908 6502 4910 6554
rect 5090 6502 5092 6554
rect 4846 6500 4852 6502
rect 4908 6500 4932 6502
rect 4988 6500 5012 6502
rect 5068 6500 5092 6502
rect 5148 6500 5154 6502
rect 4846 6491 5154 6500
rect 6794 6556 7102 6565
rect 6794 6554 6800 6556
rect 6856 6554 6880 6556
rect 6936 6554 6960 6556
rect 7016 6554 7040 6556
rect 7096 6554 7102 6556
rect 6856 6502 6858 6554
rect 7038 6502 7040 6554
rect 6794 6500 6800 6502
rect 6856 6500 6880 6502
rect 6936 6500 6960 6502
rect 7016 6500 7040 6502
rect 7096 6500 7102 6502
rect 6794 6491 7102 6500
rect 1924 6012 2232 6021
rect 1924 6010 1930 6012
rect 1986 6010 2010 6012
rect 2066 6010 2090 6012
rect 2146 6010 2170 6012
rect 2226 6010 2232 6012
rect 1986 5958 1988 6010
rect 2168 5958 2170 6010
rect 1924 5956 1930 5958
rect 1986 5956 2010 5958
rect 2066 5956 2090 5958
rect 2146 5956 2170 5958
rect 2226 5956 2232 5958
rect 1924 5947 2232 5956
rect 3872 6012 4180 6021
rect 3872 6010 3878 6012
rect 3934 6010 3958 6012
rect 4014 6010 4038 6012
rect 4094 6010 4118 6012
rect 4174 6010 4180 6012
rect 3934 5958 3936 6010
rect 4116 5958 4118 6010
rect 3872 5956 3878 5958
rect 3934 5956 3958 5958
rect 4014 5956 4038 5958
rect 4094 5956 4118 5958
rect 4174 5956 4180 5958
rect 3872 5947 4180 5956
rect 5820 6012 6128 6021
rect 5820 6010 5826 6012
rect 5882 6010 5906 6012
rect 5962 6010 5986 6012
rect 6042 6010 6066 6012
rect 6122 6010 6128 6012
rect 5882 5958 5884 6010
rect 6064 5958 6066 6010
rect 5820 5956 5826 5958
rect 5882 5956 5906 5958
rect 5962 5956 5986 5958
rect 6042 5956 6066 5958
rect 6122 5956 6128 5958
rect 5820 5947 6128 5956
rect 7484 5710 7512 7278
rect 7768 7100 8076 7109
rect 7768 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7934 7100
rect 7990 7098 8014 7100
rect 8070 7098 8076 7100
rect 7830 7046 7832 7098
rect 8012 7046 8014 7098
rect 7768 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7934 7046
rect 7990 7044 8014 7046
rect 8070 7044 8076 7046
rect 7768 7035 8076 7044
rect 8128 6866 8156 7278
rect 9692 6866 9720 9200
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 7768 6012 8076 6021
rect 7768 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7934 6012
rect 7990 6010 8014 6012
rect 8070 6010 8076 6012
rect 7830 5958 7832 6010
rect 8012 5958 8014 6010
rect 7768 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7934 5958
rect 7990 5956 8014 5958
rect 8070 5956 8076 5958
rect 7768 5947 8076 5956
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 2898 5468 3206 5477
rect 2898 5466 2904 5468
rect 2960 5466 2984 5468
rect 3040 5466 3064 5468
rect 3120 5466 3144 5468
rect 3200 5466 3206 5468
rect 2960 5414 2962 5466
rect 3142 5414 3144 5466
rect 2898 5412 2904 5414
rect 2960 5412 2984 5414
rect 3040 5412 3064 5414
rect 3120 5412 3144 5414
rect 3200 5412 3206 5414
rect 2898 5403 3206 5412
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1924 4924 2232 4933
rect 1924 4922 1930 4924
rect 1986 4922 2010 4924
rect 2066 4922 2090 4924
rect 2146 4922 2170 4924
rect 2226 4922 2232 4924
rect 1986 4870 1988 4922
rect 2168 4870 2170 4922
rect 1924 4868 1930 4870
rect 1986 4868 2010 4870
rect 2066 4868 2090 4870
rect 2146 4868 2170 4870
rect 2226 4868 2232 4870
rect 1924 4859 2232 4868
rect 3620 4826 3648 5034
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3528 4706 3556 4762
rect 3712 4706 3740 5170
rect 3528 4678 3740 4706
rect 3712 4622 3740 4678
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3804 4554 3832 5170
rect 3872 4924 4180 4933
rect 3872 4922 3878 4924
rect 3934 4922 3958 4924
rect 4014 4922 4038 4924
rect 4094 4922 4118 4924
rect 4174 4922 4180 4924
rect 3934 4870 3936 4922
rect 4116 4870 4118 4922
rect 3872 4868 3878 4870
rect 3934 4868 3958 4870
rect 4014 4868 4038 4870
rect 4094 4868 4118 4870
rect 4174 4868 4180 4870
rect 3872 4859 4180 4868
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 2898 4380 3206 4389
rect 2898 4378 2904 4380
rect 2960 4378 2984 4380
rect 3040 4378 3064 4380
rect 3120 4378 3144 4380
rect 3200 4378 3206 4380
rect 2960 4326 2962 4378
rect 3142 4326 3144 4378
rect 2898 4324 2904 4326
rect 2960 4324 2984 4326
rect 3040 4324 3064 4326
rect 3120 4324 3144 4326
rect 3200 4324 3206 4326
rect 2898 4315 3206 4324
rect 3804 4282 3832 4490
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 4080 4010 4108 4558
rect 4172 4486 4200 4762
rect 4264 4758 4292 5170
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4146 4200 4422
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 1924 3836 2232 3845
rect 1924 3834 1930 3836
rect 1986 3834 2010 3836
rect 2066 3834 2090 3836
rect 2146 3834 2170 3836
rect 2226 3834 2232 3836
rect 1986 3782 1988 3834
rect 2168 3782 2170 3834
rect 1924 3780 1930 3782
rect 1986 3780 2010 3782
rect 2066 3780 2090 3782
rect 2146 3780 2170 3782
rect 2226 3780 2232 3782
rect 1924 3771 2232 3780
rect 2898 3292 3206 3301
rect 2898 3290 2904 3292
rect 2960 3290 2984 3292
rect 3040 3290 3064 3292
rect 3120 3290 3144 3292
rect 3200 3290 3206 3292
rect 2960 3238 2962 3290
rect 3142 3238 3144 3290
rect 2898 3236 2904 3238
rect 2960 3236 2984 3238
rect 3040 3236 3064 3238
rect 3120 3236 3144 3238
rect 3200 3236 3206 3238
rect 2898 3227 3206 3236
rect 3712 2990 3740 3878
rect 3804 3058 3832 3946
rect 3872 3836 4180 3845
rect 3872 3834 3878 3836
rect 3934 3834 3958 3836
rect 4014 3834 4038 3836
rect 4094 3834 4118 3836
rect 4174 3834 4180 3836
rect 3934 3782 3936 3834
rect 4116 3782 4118 3834
rect 3872 3780 3878 3782
rect 3934 3780 3958 3782
rect 4014 3780 4038 3782
rect 4094 3780 4118 3782
rect 4174 3780 4180 3782
rect 3872 3771 4180 3780
rect 4356 3534 4384 5646
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4632 5370 4660 5578
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 4846 5468 5154 5477
rect 4846 5466 4852 5468
rect 4908 5466 4932 5468
rect 4988 5466 5012 5468
rect 5068 5466 5092 5468
rect 5148 5466 5154 5468
rect 4908 5414 4910 5466
rect 5090 5414 5092 5466
rect 4846 5412 4852 5414
rect 4908 5412 4932 5414
rect 4988 5412 5012 5414
rect 5068 5412 5092 5414
rect 5148 5412 5154 5414
rect 4846 5403 5154 5412
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4724 4826 4752 5238
rect 5820 4924 6128 4933
rect 5820 4922 5826 4924
rect 5882 4922 5906 4924
rect 5962 4922 5986 4924
rect 6042 4922 6066 4924
rect 6122 4922 6128 4924
rect 5882 4870 5884 4922
rect 6064 4870 6066 4922
rect 5820 4868 5826 4870
rect 5882 4868 5906 4870
rect 5962 4868 5986 4870
rect 6042 4868 6066 4870
rect 6122 4868 6128 4870
rect 5820 4859 6128 4868
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4632 4146 4660 4626
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 4846 4380 5154 4389
rect 4846 4378 4852 4380
rect 4908 4378 4932 4380
rect 4988 4378 5012 4380
rect 5068 4378 5092 4380
rect 5148 4378 5154 4380
rect 4908 4326 4910 4378
rect 5090 4326 5092 4378
rect 4846 4324 4852 4326
rect 4908 4324 4932 4326
rect 4988 4324 5012 4326
rect 5068 4324 5092 4326
rect 5148 4324 5154 4326
rect 4846 4315 5154 4324
rect 5552 4282 5580 4558
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4632 3738 4660 4082
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 5736 3534 5764 3878
rect 5820 3836 6128 3845
rect 5820 3834 5826 3836
rect 5882 3834 5906 3836
rect 5962 3834 5986 3836
rect 6042 3834 6066 3836
rect 6122 3834 6128 3836
rect 5882 3782 5884 3834
rect 6064 3782 6066 3834
rect 5820 3780 5826 3782
rect 5882 3780 5906 3782
rect 5962 3780 5986 3782
rect 6042 3780 6066 3782
rect 6122 3780 6128 3782
rect 5820 3771 6128 3780
rect 6196 3602 6224 4558
rect 6564 3942 6592 5510
rect 6794 5468 7102 5477
rect 6794 5466 6800 5468
rect 6856 5466 6880 5468
rect 6936 5466 6960 5468
rect 7016 5466 7040 5468
rect 7096 5466 7102 5468
rect 6856 5414 6858 5466
rect 7038 5414 7040 5466
rect 6794 5412 6800 5414
rect 6856 5412 6880 5414
rect 6936 5412 6960 5414
rect 7016 5412 7040 5414
rect 7096 5412 7102 5414
rect 6794 5403 7102 5412
rect 7484 5234 7512 5646
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 5114 7512 5170
rect 7392 5086 7512 5114
rect 6794 4380 7102 4389
rect 6794 4378 6800 4380
rect 6856 4378 6880 4380
rect 6936 4378 6960 4380
rect 7016 4378 7040 4380
rect 7096 4378 7102 4380
rect 6856 4326 6858 4378
rect 7038 4326 7040 4378
rect 6794 4324 6800 4326
rect 6856 4324 6880 4326
rect 6936 4324 6960 4326
rect 7016 4324 7040 4326
rect 7096 4324 7102 4326
rect 6794 4315 7102 4324
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4172 2990 4200 3402
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 1924 2748 2232 2757
rect 1924 2746 1930 2748
rect 1986 2746 2010 2748
rect 2066 2746 2090 2748
rect 2146 2746 2170 2748
rect 2226 2746 2232 2748
rect 1986 2694 1988 2746
rect 2168 2694 2170 2746
rect 1924 2692 1930 2694
rect 1986 2692 2010 2694
rect 2066 2692 2090 2694
rect 2146 2692 2170 2694
rect 2226 2692 2232 2694
rect 1924 2683 2232 2692
rect 3872 2748 4180 2757
rect 3872 2746 3878 2748
rect 3934 2746 3958 2748
rect 4014 2746 4038 2748
rect 4094 2746 4118 2748
rect 4174 2746 4180 2748
rect 3934 2694 3936 2746
rect 4116 2694 4118 2746
rect 3872 2692 3878 2694
rect 3934 2692 3958 2694
rect 4014 2692 4038 2694
rect 4094 2692 4118 2694
rect 4174 2692 4180 2694
rect 3872 2683 4180 2692
rect 4356 2650 4384 3470
rect 4846 3292 5154 3301
rect 4846 3290 4852 3292
rect 4908 3290 4932 3292
rect 4988 3290 5012 3292
rect 5068 3290 5092 3292
rect 5148 3290 5154 3292
rect 4908 3238 4910 3290
rect 5090 3238 5092 3290
rect 4846 3236 4852 3238
rect 4908 3236 4932 3238
rect 4988 3236 5012 3238
rect 5068 3236 5092 3238
rect 5148 3236 5154 3238
rect 4846 3227 5154 3236
rect 6656 3074 6684 4150
rect 7392 4146 7420 5086
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4554 7512 4966
rect 7768 4924 8076 4933
rect 7768 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7934 4924
rect 7990 4922 8014 4924
rect 8070 4922 8076 4924
rect 7830 4870 7832 4922
rect 8012 4870 8014 4922
rect 7768 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7934 4870
rect 7990 4868 8014 4870
rect 8070 4868 8076 4870
rect 7768 4859 8076 4868
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6932 3738 6960 3946
rect 7768 3836 8076 3845
rect 7768 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7934 3836
rect 7990 3834 8014 3836
rect 8070 3834 8076 3836
rect 7830 3782 7832 3834
rect 8012 3782 8014 3834
rect 7768 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7934 3782
rect 7990 3780 8014 3782
rect 8070 3780 8076 3782
rect 7768 3771 8076 3780
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6794 3292 7102 3301
rect 6794 3290 6800 3292
rect 6856 3290 6880 3292
rect 6936 3290 6960 3292
rect 7016 3290 7040 3292
rect 7096 3290 7102 3292
rect 6856 3238 6858 3290
rect 7038 3238 7040 3290
rect 6794 3236 6800 3238
rect 6856 3236 6880 3238
rect 6936 3236 6960 3238
rect 7016 3236 7040 3238
rect 7096 3236 7102 3238
rect 6794 3227 7102 3236
rect 6656 3046 6960 3074
rect 5820 2748 6128 2757
rect 5820 2746 5826 2748
rect 5882 2746 5906 2748
rect 5962 2746 5986 2748
rect 6042 2746 6066 2748
rect 6122 2746 6128 2748
rect 5882 2694 5884 2746
rect 6064 2694 6066 2746
rect 5820 2692 5826 2694
rect 5882 2692 5906 2694
rect 5962 2692 5986 2694
rect 6042 2692 6066 2694
rect 6122 2692 6128 2694
rect 5820 2683 6128 2692
rect 6932 2650 6960 3046
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 7768 2748 8076 2757
rect 7768 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7934 2748
rect 7990 2746 8014 2748
rect 8070 2746 8076 2748
rect 7830 2694 7832 2746
rect 8012 2694 8014 2746
rect 7768 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7934 2694
rect 7990 2692 8014 2694
rect 8070 2692 8076 2694
rect 7768 2683 8076 2692
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 8128 2446 8156 2790
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 32 800 60 2382
rect 2898 2204 3206 2213
rect 2898 2202 2904 2204
rect 2960 2202 2984 2204
rect 3040 2202 3064 2204
rect 3120 2202 3144 2204
rect 3200 2202 3206 2204
rect 2960 2150 2962 2202
rect 3142 2150 3144 2202
rect 2898 2148 2904 2150
rect 2960 2148 2984 2150
rect 3040 2148 3064 2150
rect 3120 2148 3144 2150
rect 3200 2148 3206 2150
rect 2898 2139 3206 2148
rect 4846 2204 5154 2213
rect 4846 2202 4852 2204
rect 4908 2202 4932 2204
rect 4988 2202 5012 2204
rect 5068 2202 5092 2204
rect 5148 2202 5154 2204
rect 4908 2150 4910 2202
rect 5090 2150 5092 2202
rect 4846 2148 4852 2150
rect 4908 2148 4932 2150
rect 4988 2148 5012 2150
rect 5068 2148 5092 2150
rect 5148 2148 5154 2150
rect 4846 2139 5154 2148
rect 6794 2204 7102 2213
rect 6794 2202 6800 2204
rect 6856 2202 6880 2204
rect 6936 2202 6960 2204
rect 7016 2202 7040 2204
rect 7096 2202 7102 2204
rect 6856 2150 6858 2202
rect 7038 2150 7040 2202
rect 6794 2148 6800 2150
rect 6856 2148 6880 2150
rect 6936 2148 6960 2150
rect 7016 2148 7040 2150
rect 7096 2148 7102 2150
rect 6794 2139 7102 2148
rect 9692 800 9720 2790
rect 18 0 74 800
rect 9678 0 9734 800
<< via2 >>
rect 2904 7642 2960 7644
rect 2984 7642 3040 7644
rect 3064 7642 3120 7644
rect 3144 7642 3200 7644
rect 2904 7590 2950 7642
rect 2950 7590 2960 7642
rect 2984 7590 3014 7642
rect 3014 7590 3026 7642
rect 3026 7590 3040 7642
rect 3064 7590 3078 7642
rect 3078 7590 3090 7642
rect 3090 7590 3120 7642
rect 3144 7590 3154 7642
rect 3154 7590 3200 7642
rect 2904 7588 2960 7590
rect 2984 7588 3040 7590
rect 3064 7588 3120 7590
rect 3144 7588 3200 7590
rect 4852 7642 4908 7644
rect 4932 7642 4988 7644
rect 5012 7642 5068 7644
rect 5092 7642 5148 7644
rect 4852 7590 4898 7642
rect 4898 7590 4908 7642
rect 4932 7590 4962 7642
rect 4962 7590 4974 7642
rect 4974 7590 4988 7642
rect 5012 7590 5026 7642
rect 5026 7590 5038 7642
rect 5038 7590 5068 7642
rect 5092 7590 5102 7642
rect 5102 7590 5148 7642
rect 4852 7588 4908 7590
rect 4932 7588 4988 7590
rect 5012 7588 5068 7590
rect 5092 7588 5148 7590
rect 6800 7642 6856 7644
rect 6880 7642 6936 7644
rect 6960 7642 7016 7644
rect 7040 7642 7096 7644
rect 6800 7590 6846 7642
rect 6846 7590 6856 7642
rect 6880 7590 6910 7642
rect 6910 7590 6922 7642
rect 6922 7590 6936 7642
rect 6960 7590 6974 7642
rect 6974 7590 6986 7642
rect 6986 7590 7016 7642
rect 7040 7590 7050 7642
rect 7050 7590 7096 7642
rect 6800 7588 6856 7590
rect 6880 7588 6936 7590
rect 6960 7588 7016 7590
rect 7040 7588 7096 7590
rect 1930 7098 1986 7100
rect 2010 7098 2066 7100
rect 2090 7098 2146 7100
rect 2170 7098 2226 7100
rect 1930 7046 1976 7098
rect 1976 7046 1986 7098
rect 2010 7046 2040 7098
rect 2040 7046 2052 7098
rect 2052 7046 2066 7098
rect 2090 7046 2104 7098
rect 2104 7046 2116 7098
rect 2116 7046 2146 7098
rect 2170 7046 2180 7098
rect 2180 7046 2226 7098
rect 1930 7044 1986 7046
rect 2010 7044 2066 7046
rect 2090 7044 2146 7046
rect 2170 7044 2226 7046
rect 3878 7098 3934 7100
rect 3958 7098 4014 7100
rect 4038 7098 4094 7100
rect 4118 7098 4174 7100
rect 3878 7046 3924 7098
rect 3924 7046 3934 7098
rect 3958 7046 3988 7098
rect 3988 7046 4000 7098
rect 4000 7046 4014 7098
rect 4038 7046 4052 7098
rect 4052 7046 4064 7098
rect 4064 7046 4094 7098
rect 4118 7046 4128 7098
rect 4128 7046 4174 7098
rect 3878 7044 3934 7046
rect 3958 7044 4014 7046
rect 4038 7044 4094 7046
rect 4118 7044 4174 7046
rect 5826 7098 5882 7100
rect 5906 7098 5962 7100
rect 5986 7098 6042 7100
rect 6066 7098 6122 7100
rect 5826 7046 5872 7098
rect 5872 7046 5882 7098
rect 5906 7046 5936 7098
rect 5936 7046 5948 7098
rect 5948 7046 5962 7098
rect 5986 7046 6000 7098
rect 6000 7046 6012 7098
rect 6012 7046 6042 7098
rect 6066 7046 6076 7098
rect 6076 7046 6122 7098
rect 5826 7044 5882 7046
rect 5906 7044 5962 7046
rect 5986 7044 6042 7046
rect 6066 7044 6122 7046
rect 2904 6554 2960 6556
rect 2984 6554 3040 6556
rect 3064 6554 3120 6556
rect 3144 6554 3200 6556
rect 2904 6502 2950 6554
rect 2950 6502 2960 6554
rect 2984 6502 3014 6554
rect 3014 6502 3026 6554
rect 3026 6502 3040 6554
rect 3064 6502 3078 6554
rect 3078 6502 3090 6554
rect 3090 6502 3120 6554
rect 3144 6502 3154 6554
rect 3154 6502 3200 6554
rect 2904 6500 2960 6502
rect 2984 6500 3040 6502
rect 3064 6500 3120 6502
rect 3144 6500 3200 6502
rect 4852 6554 4908 6556
rect 4932 6554 4988 6556
rect 5012 6554 5068 6556
rect 5092 6554 5148 6556
rect 4852 6502 4898 6554
rect 4898 6502 4908 6554
rect 4932 6502 4962 6554
rect 4962 6502 4974 6554
rect 4974 6502 4988 6554
rect 5012 6502 5026 6554
rect 5026 6502 5038 6554
rect 5038 6502 5068 6554
rect 5092 6502 5102 6554
rect 5102 6502 5148 6554
rect 4852 6500 4908 6502
rect 4932 6500 4988 6502
rect 5012 6500 5068 6502
rect 5092 6500 5148 6502
rect 6800 6554 6856 6556
rect 6880 6554 6936 6556
rect 6960 6554 7016 6556
rect 7040 6554 7096 6556
rect 6800 6502 6846 6554
rect 6846 6502 6856 6554
rect 6880 6502 6910 6554
rect 6910 6502 6922 6554
rect 6922 6502 6936 6554
rect 6960 6502 6974 6554
rect 6974 6502 6986 6554
rect 6986 6502 7016 6554
rect 7040 6502 7050 6554
rect 7050 6502 7096 6554
rect 6800 6500 6856 6502
rect 6880 6500 6936 6502
rect 6960 6500 7016 6502
rect 7040 6500 7096 6502
rect 1930 6010 1986 6012
rect 2010 6010 2066 6012
rect 2090 6010 2146 6012
rect 2170 6010 2226 6012
rect 1930 5958 1976 6010
rect 1976 5958 1986 6010
rect 2010 5958 2040 6010
rect 2040 5958 2052 6010
rect 2052 5958 2066 6010
rect 2090 5958 2104 6010
rect 2104 5958 2116 6010
rect 2116 5958 2146 6010
rect 2170 5958 2180 6010
rect 2180 5958 2226 6010
rect 1930 5956 1986 5958
rect 2010 5956 2066 5958
rect 2090 5956 2146 5958
rect 2170 5956 2226 5958
rect 3878 6010 3934 6012
rect 3958 6010 4014 6012
rect 4038 6010 4094 6012
rect 4118 6010 4174 6012
rect 3878 5958 3924 6010
rect 3924 5958 3934 6010
rect 3958 5958 3988 6010
rect 3988 5958 4000 6010
rect 4000 5958 4014 6010
rect 4038 5958 4052 6010
rect 4052 5958 4064 6010
rect 4064 5958 4094 6010
rect 4118 5958 4128 6010
rect 4128 5958 4174 6010
rect 3878 5956 3934 5958
rect 3958 5956 4014 5958
rect 4038 5956 4094 5958
rect 4118 5956 4174 5958
rect 5826 6010 5882 6012
rect 5906 6010 5962 6012
rect 5986 6010 6042 6012
rect 6066 6010 6122 6012
rect 5826 5958 5872 6010
rect 5872 5958 5882 6010
rect 5906 5958 5936 6010
rect 5936 5958 5948 6010
rect 5948 5958 5962 6010
rect 5986 5958 6000 6010
rect 6000 5958 6012 6010
rect 6012 5958 6042 6010
rect 6066 5958 6076 6010
rect 6076 5958 6122 6010
rect 5826 5956 5882 5958
rect 5906 5956 5962 5958
rect 5986 5956 6042 5958
rect 6066 5956 6122 5958
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7934 7098 7990 7100
rect 8014 7098 8070 7100
rect 7774 7046 7820 7098
rect 7820 7046 7830 7098
rect 7854 7046 7884 7098
rect 7884 7046 7896 7098
rect 7896 7046 7910 7098
rect 7934 7046 7948 7098
rect 7948 7046 7960 7098
rect 7960 7046 7990 7098
rect 8014 7046 8024 7098
rect 8024 7046 8070 7098
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7934 7044 7990 7046
rect 8014 7044 8070 7046
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7934 6010 7990 6012
rect 8014 6010 8070 6012
rect 7774 5958 7820 6010
rect 7820 5958 7830 6010
rect 7854 5958 7884 6010
rect 7884 5958 7896 6010
rect 7896 5958 7910 6010
rect 7934 5958 7948 6010
rect 7948 5958 7960 6010
rect 7960 5958 7990 6010
rect 8014 5958 8024 6010
rect 8024 5958 8070 6010
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 7934 5956 7990 5958
rect 8014 5956 8070 5958
rect 2904 5466 2960 5468
rect 2984 5466 3040 5468
rect 3064 5466 3120 5468
rect 3144 5466 3200 5468
rect 2904 5414 2950 5466
rect 2950 5414 2960 5466
rect 2984 5414 3014 5466
rect 3014 5414 3026 5466
rect 3026 5414 3040 5466
rect 3064 5414 3078 5466
rect 3078 5414 3090 5466
rect 3090 5414 3120 5466
rect 3144 5414 3154 5466
rect 3154 5414 3200 5466
rect 2904 5412 2960 5414
rect 2984 5412 3040 5414
rect 3064 5412 3120 5414
rect 3144 5412 3200 5414
rect 1930 4922 1986 4924
rect 2010 4922 2066 4924
rect 2090 4922 2146 4924
rect 2170 4922 2226 4924
rect 1930 4870 1976 4922
rect 1976 4870 1986 4922
rect 2010 4870 2040 4922
rect 2040 4870 2052 4922
rect 2052 4870 2066 4922
rect 2090 4870 2104 4922
rect 2104 4870 2116 4922
rect 2116 4870 2146 4922
rect 2170 4870 2180 4922
rect 2180 4870 2226 4922
rect 1930 4868 1986 4870
rect 2010 4868 2066 4870
rect 2090 4868 2146 4870
rect 2170 4868 2226 4870
rect 3878 4922 3934 4924
rect 3958 4922 4014 4924
rect 4038 4922 4094 4924
rect 4118 4922 4174 4924
rect 3878 4870 3924 4922
rect 3924 4870 3934 4922
rect 3958 4870 3988 4922
rect 3988 4870 4000 4922
rect 4000 4870 4014 4922
rect 4038 4870 4052 4922
rect 4052 4870 4064 4922
rect 4064 4870 4094 4922
rect 4118 4870 4128 4922
rect 4128 4870 4174 4922
rect 3878 4868 3934 4870
rect 3958 4868 4014 4870
rect 4038 4868 4094 4870
rect 4118 4868 4174 4870
rect 2904 4378 2960 4380
rect 2984 4378 3040 4380
rect 3064 4378 3120 4380
rect 3144 4378 3200 4380
rect 2904 4326 2950 4378
rect 2950 4326 2960 4378
rect 2984 4326 3014 4378
rect 3014 4326 3026 4378
rect 3026 4326 3040 4378
rect 3064 4326 3078 4378
rect 3078 4326 3090 4378
rect 3090 4326 3120 4378
rect 3144 4326 3154 4378
rect 3154 4326 3200 4378
rect 2904 4324 2960 4326
rect 2984 4324 3040 4326
rect 3064 4324 3120 4326
rect 3144 4324 3200 4326
rect 1930 3834 1986 3836
rect 2010 3834 2066 3836
rect 2090 3834 2146 3836
rect 2170 3834 2226 3836
rect 1930 3782 1976 3834
rect 1976 3782 1986 3834
rect 2010 3782 2040 3834
rect 2040 3782 2052 3834
rect 2052 3782 2066 3834
rect 2090 3782 2104 3834
rect 2104 3782 2116 3834
rect 2116 3782 2146 3834
rect 2170 3782 2180 3834
rect 2180 3782 2226 3834
rect 1930 3780 1986 3782
rect 2010 3780 2066 3782
rect 2090 3780 2146 3782
rect 2170 3780 2226 3782
rect 2904 3290 2960 3292
rect 2984 3290 3040 3292
rect 3064 3290 3120 3292
rect 3144 3290 3200 3292
rect 2904 3238 2950 3290
rect 2950 3238 2960 3290
rect 2984 3238 3014 3290
rect 3014 3238 3026 3290
rect 3026 3238 3040 3290
rect 3064 3238 3078 3290
rect 3078 3238 3090 3290
rect 3090 3238 3120 3290
rect 3144 3238 3154 3290
rect 3154 3238 3200 3290
rect 2904 3236 2960 3238
rect 2984 3236 3040 3238
rect 3064 3236 3120 3238
rect 3144 3236 3200 3238
rect 3878 3834 3934 3836
rect 3958 3834 4014 3836
rect 4038 3834 4094 3836
rect 4118 3834 4174 3836
rect 3878 3782 3924 3834
rect 3924 3782 3934 3834
rect 3958 3782 3988 3834
rect 3988 3782 4000 3834
rect 4000 3782 4014 3834
rect 4038 3782 4052 3834
rect 4052 3782 4064 3834
rect 4064 3782 4094 3834
rect 4118 3782 4128 3834
rect 4128 3782 4174 3834
rect 3878 3780 3934 3782
rect 3958 3780 4014 3782
rect 4038 3780 4094 3782
rect 4118 3780 4174 3782
rect 4852 5466 4908 5468
rect 4932 5466 4988 5468
rect 5012 5466 5068 5468
rect 5092 5466 5148 5468
rect 4852 5414 4898 5466
rect 4898 5414 4908 5466
rect 4932 5414 4962 5466
rect 4962 5414 4974 5466
rect 4974 5414 4988 5466
rect 5012 5414 5026 5466
rect 5026 5414 5038 5466
rect 5038 5414 5068 5466
rect 5092 5414 5102 5466
rect 5102 5414 5148 5466
rect 4852 5412 4908 5414
rect 4932 5412 4988 5414
rect 5012 5412 5068 5414
rect 5092 5412 5148 5414
rect 5826 4922 5882 4924
rect 5906 4922 5962 4924
rect 5986 4922 6042 4924
rect 6066 4922 6122 4924
rect 5826 4870 5872 4922
rect 5872 4870 5882 4922
rect 5906 4870 5936 4922
rect 5936 4870 5948 4922
rect 5948 4870 5962 4922
rect 5986 4870 6000 4922
rect 6000 4870 6012 4922
rect 6012 4870 6042 4922
rect 6066 4870 6076 4922
rect 6076 4870 6122 4922
rect 5826 4868 5882 4870
rect 5906 4868 5962 4870
rect 5986 4868 6042 4870
rect 6066 4868 6122 4870
rect 4852 4378 4908 4380
rect 4932 4378 4988 4380
rect 5012 4378 5068 4380
rect 5092 4378 5148 4380
rect 4852 4326 4898 4378
rect 4898 4326 4908 4378
rect 4932 4326 4962 4378
rect 4962 4326 4974 4378
rect 4974 4326 4988 4378
rect 5012 4326 5026 4378
rect 5026 4326 5038 4378
rect 5038 4326 5068 4378
rect 5092 4326 5102 4378
rect 5102 4326 5148 4378
rect 4852 4324 4908 4326
rect 4932 4324 4988 4326
rect 5012 4324 5068 4326
rect 5092 4324 5148 4326
rect 5826 3834 5882 3836
rect 5906 3834 5962 3836
rect 5986 3834 6042 3836
rect 6066 3834 6122 3836
rect 5826 3782 5872 3834
rect 5872 3782 5882 3834
rect 5906 3782 5936 3834
rect 5936 3782 5948 3834
rect 5948 3782 5962 3834
rect 5986 3782 6000 3834
rect 6000 3782 6012 3834
rect 6012 3782 6042 3834
rect 6066 3782 6076 3834
rect 6076 3782 6122 3834
rect 5826 3780 5882 3782
rect 5906 3780 5962 3782
rect 5986 3780 6042 3782
rect 6066 3780 6122 3782
rect 6800 5466 6856 5468
rect 6880 5466 6936 5468
rect 6960 5466 7016 5468
rect 7040 5466 7096 5468
rect 6800 5414 6846 5466
rect 6846 5414 6856 5466
rect 6880 5414 6910 5466
rect 6910 5414 6922 5466
rect 6922 5414 6936 5466
rect 6960 5414 6974 5466
rect 6974 5414 6986 5466
rect 6986 5414 7016 5466
rect 7040 5414 7050 5466
rect 7050 5414 7096 5466
rect 6800 5412 6856 5414
rect 6880 5412 6936 5414
rect 6960 5412 7016 5414
rect 7040 5412 7096 5414
rect 6800 4378 6856 4380
rect 6880 4378 6936 4380
rect 6960 4378 7016 4380
rect 7040 4378 7096 4380
rect 6800 4326 6846 4378
rect 6846 4326 6856 4378
rect 6880 4326 6910 4378
rect 6910 4326 6922 4378
rect 6922 4326 6936 4378
rect 6960 4326 6974 4378
rect 6974 4326 6986 4378
rect 6986 4326 7016 4378
rect 7040 4326 7050 4378
rect 7050 4326 7096 4378
rect 6800 4324 6856 4326
rect 6880 4324 6936 4326
rect 6960 4324 7016 4326
rect 7040 4324 7096 4326
rect 1930 2746 1986 2748
rect 2010 2746 2066 2748
rect 2090 2746 2146 2748
rect 2170 2746 2226 2748
rect 1930 2694 1976 2746
rect 1976 2694 1986 2746
rect 2010 2694 2040 2746
rect 2040 2694 2052 2746
rect 2052 2694 2066 2746
rect 2090 2694 2104 2746
rect 2104 2694 2116 2746
rect 2116 2694 2146 2746
rect 2170 2694 2180 2746
rect 2180 2694 2226 2746
rect 1930 2692 1986 2694
rect 2010 2692 2066 2694
rect 2090 2692 2146 2694
rect 2170 2692 2226 2694
rect 3878 2746 3934 2748
rect 3958 2746 4014 2748
rect 4038 2746 4094 2748
rect 4118 2746 4174 2748
rect 3878 2694 3924 2746
rect 3924 2694 3934 2746
rect 3958 2694 3988 2746
rect 3988 2694 4000 2746
rect 4000 2694 4014 2746
rect 4038 2694 4052 2746
rect 4052 2694 4064 2746
rect 4064 2694 4094 2746
rect 4118 2694 4128 2746
rect 4128 2694 4174 2746
rect 3878 2692 3934 2694
rect 3958 2692 4014 2694
rect 4038 2692 4094 2694
rect 4118 2692 4174 2694
rect 4852 3290 4908 3292
rect 4932 3290 4988 3292
rect 5012 3290 5068 3292
rect 5092 3290 5148 3292
rect 4852 3238 4898 3290
rect 4898 3238 4908 3290
rect 4932 3238 4962 3290
rect 4962 3238 4974 3290
rect 4974 3238 4988 3290
rect 5012 3238 5026 3290
rect 5026 3238 5038 3290
rect 5038 3238 5068 3290
rect 5092 3238 5102 3290
rect 5102 3238 5148 3290
rect 4852 3236 4908 3238
rect 4932 3236 4988 3238
rect 5012 3236 5068 3238
rect 5092 3236 5148 3238
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7934 4922 7990 4924
rect 8014 4922 8070 4924
rect 7774 4870 7820 4922
rect 7820 4870 7830 4922
rect 7854 4870 7884 4922
rect 7884 4870 7896 4922
rect 7896 4870 7910 4922
rect 7934 4870 7948 4922
rect 7948 4870 7960 4922
rect 7960 4870 7990 4922
rect 8014 4870 8024 4922
rect 8024 4870 8070 4922
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 7934 4868 7990 4870
rect 8014 4868 8070 4870
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7934 3834 7990 3836
rect 8014 3834 8070 3836
rect 7774 3782 7820 3834
rect 7820 3782 7830 3834
rect 7854 3782 7884 3834
rect 7884 3782 7896 3834
rect 7896 3782 7910 3834
rect 7934 3782 7948 3834
rect 7948 3782 7960 3834
rect 7960 3782 7990 3834
rect 8014 3782 8024 3834
rect 8024 3782 8070 3834
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 7934 3780 7990 3782
rect 8014 3780 8070 3782
rect 6800 3290 6856 3292
rect 6880 3290 6936 3292
rect 6960 3290 7016 3292
rect 7040 3290 7096 3292
rect 6800 3238 6846 3290
rect 6846 3238 6856 3290
rect 6880 3238 6910 3290
rect 6910 3238 6922 3290
rect 6922 3238 6936 3290
rect 6960 3238 6974 3290
rect 6974 3238 6986 3290
rect 6986 3238 7016 3290
rect 7040 3238 7050 3290
rect 7050 3238 7096 3290
rect 6800 3236 6856 3238
rect 6880 3236 6936 3238
rect 6960 3236 7016 3238
rect 7040 3236 7096 3238
rect 5826 2746 5882 2748
rect 5906 2746 5962 2748
rect 5986 2746 6042 2748
rect 6066 2746 6122 2748
rect 5826 2694 5872 2746
rect 5872 2694 5882 2746
rect 5906 2694 5936 2746
rect 5936 2694 5948 2746
rect 5948 2694 5962 2746
rect 5986 2694 6000 2746
rect 6000 2694 6012 2746
rect 6012 2694 6042 2746
rect 6066 2694 6076 2746
rect 6076 2694 6122 2746
rect 5826 2692 5882 2694
rect 5906 2692 5962 2694
rect 5986 2692 6042 2694
rect 6066 2692 6122 2694
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7934 2746 7990 2748
rect 8014 2746 8070 2748
rect 7774 2694 7820 2746
rect 7820 2694 7830 2746
rect 7854 2694 7884 2746
rect 7884 2694 7896 2746
rect 7896 2694 7910 2746
rect 7934 2694 7948 2746
rect 7948 2694 7960 2746
rect 7960 2694 7990 2746
rect 8014 2694 8024 2746
rect 8024 2694 8070 2746
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 7934 2692 7990 2694
rect 8014 2692 8070 2694
rect 2904 2202 2960 2204
rect 2984 2202 3040 2204
rect 3064 2202 3120 2204
rect 3144 2202 3200 2204
rect 2904 2150 2950 2202
rect 2950 2150 2960 2202
rect 2984 2150 3014 2202
rect 3014 2150 3026 2202
rect 3026 2150 3040 2202
rect 3064 2150 3078 2202
rect 3078 2150 3090 2202
rect 3090 2150 3120 2202
rect 3144 2150 3154 2202
rect 3154 2150 3200 2202
rect 2904 2148 2960 2150
rect 2984 2148 3040 2150
rect 3064 2148 3120 2150
rect 3144 2148 3200 2150
rect 4852 2202 4908 2204
rect 4932 2202 4988 2204
rect 5012 2202 5068 2204
rect 5092 2202 5148 2204
rect 4852 2150 4898 2202
rect 4898 2150 4908 2202
rect 4932 2150 4962 2202
rect 4962 2150 4974 2202
rect 4974 2150 4988 2202
rect 5012 2150 5026 2202
rect 5026 2150 5038 2202
rect 5038 2150 5068 2202
rect 5092 2150 5102 2202
rect 5102 2150 5148 2202
rect 4852 2148 4908 2150
rect 4932 2148 4988 2150
rect 5012 2148 5068 2150
rect 5092 2148 5148 2150
rect 6800 2202 6856 2204
rect 6880 2202 6936 2204
rect 6960 2202 7016 2204
rect 7040 2202 7096 2204
rect 6800 2150 6846 2202
rect 6846 2150 6856 2202
rect 6880 2150 6910 2202
rect 6910 2150 6922 2202
rect 6922 2150 6936 2202
rect 6960 2150 6974 2202
rect 6974 2150 6986 2202
rect 6986 2150 7016 2202
rect 7040 2150 7050 2202
rect 7050 2150 7096 2202
rect 6800 2148 6856 2150
rect 6880 2148 6936 2150
rect 6960 2148 7016 2150
rect 7040 2148 7096 2150
<< metal3 >>
rect 2894 7648 3210 7649
rect 2894 7584 2900 7648
rect 2964 7584 2980 7648
rect 3044 7584 3060 7648
rect 3124 7584 3140 7648
rect 3204 7584 3210 7648
rect 2894 7583 3210 7584
rect 4842 7648 5158 7649
rect 4842 7584 4848 7648
rect 4912 7584 4928 7648
rect 4992 7584 5008 7648
rect 5072 7584 5088 7648
rect 5152 7584 5158 7648
rect 4842 7583 5158 7584
rect 6790 7648 7106 7649
rect 6790 7584 6796 7648
rect 6860 7584 6876 7648
rect 6940 7584 6956 7648
rect 7020 7584 7036 7648
rect 7100 7584 7106 7648
rect 6790 7583 7106 7584
rect 1920 7104 2236 7105
rect 1920 7040 1926 7104
rect 1990 7040 2006 7104
rect 2070 7040 2086 7104
rect 2150 7040 2166 7104
rect 2230 7040 2236 7104
rect 1920 7039 2236 7040
rect 3868 7104 4184 7105
rect 3868 7040 3874 7104
rect 3938 7040 3954 7104
rect 4018 7040 4034 7104
rect 4098 7040 4114 7104
rect 4178 7040 4184 7104
rect 3868 7039 4184 7040
rect 5816 7104 6132 7105
rect 5816 7040 5822 7104
rect 5886 7040 5902 7104
rect 5966 7040 5982 7104
rect 6046 7040 6062 7104
rect 6126 7040 6132 7104
rect 5816 7039 6132 7040
rect 7764 7104 8080 7105
rect 7764 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7930 7104
rect 7994 7040 8010 7104
rect 8074 7040 8080 7104
rect 7764 7039 8080 7040
rect 2894 6560 3210 6561
rect 2894 6496 2900 6560
rect 2964 6496 2980 6560
rect 3044 6496 3060 6560
rect 3124 6496 3140 6560
rect 3204 6496 3210 6560
rect 2894 6495 3210 6496
rect 4842 6560 5158 6561
rect 4842 6496 4848 6560
rect 4912 6496 4928 6560
rect 4992 6496 5008 6560
rect 5072 6496 5088 6560
rect 5152 6496 5158 6560
rect 4842 6495 5158 6496
rect 6790 6560 7106 6561
rect 6790 6496 6796 6560
rect 6860 6496 6876 6560
rect 6940 6496 6956 6560
rect 7020 6496 7036 6560
rect 7100 6496 7106 6560
rect 6790 6495 7106 6496
rect 1920 6016 2236 6017
rect 1920 5952 1926 6016
rect 1990 5952 2006 6016
rect 2070 5952 2086 6016
rect 2150 5952 2166 6016
rect 2230 5952 2236 6016
rect 1920 5951 2236 5952
rect 3868 6016 4184 6017
rect 3868 5952 3874 6016
rect 3938 5952 3954 6016
rect 4018 5952 4034 6016
rect 4098 5952 4114 6016
rect 4178 5952 4184 6016
rect 3868 5951 4184 5952
rect 5816 6016 6132 6017
rect 5816 5952 5822 6016
rect 5886 5952 5902 6016
rect 5966 5952 5982 6016
rect 6046 5952 6062 6016
rect 6126 5952 6132 6016
rect 5816 5951 6132 5952
rect 7764 6016 8080 6017
rect 7764 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7930 6016
rect 7994 5952 8010 6016
rect 8074 5952 8080 6016
rect 7764 5951 8080 5952
rect 2894 5472 3210 5473
rect 2894 5408 2900 5472
rect 2964 5408 2980 5472
rect 3044 5408 3060 5472
rect 3124 5408 3140 5472
rect 3204 5408 3210 5472
rect 2894 5407 3210 5408
rect 4842 5472 5158 5473
rect 4842 5408 4848 5472
rect 4912 5408 4928 5472
rect 4992 5408 5008 5472
rect 5072 5408 5088 5472
rect 5152 5408 5158 5472
rect 4842 5407 5158 5408
rect 6790 5472 7106 5473
rect 6790 5408 6796 5472
rect 6860 5408 6876 5472
rect 6940 5408 6956 5472
rect 7020 5408 7036 5472
rect 7100 5408 7106 5472
rect 6790 5407 7106 5408
rect 1920 4928 2236 4929
rect 1920 4864 1926 4928
rect 1990 4864 2006 4928
rect 2070 4864 2086 4928
rect 2150 4864 2166 4928
rect 2230 4864 2236 4928
rect 1920 4863 2236 4864
rect 3868 4928 4184 4929
rect 3868 4864 3874 4928
rect 3938 4864 3954 4928
rect 4018 4864 4034 4928
rect 4098 4864 4114 4928
rect 4178 4864 4184 4928
rect 3868 4863 4184 4864
rect 5816 4928 6132 4929
rect 5816 4864 5822 4928
rect 5886 4864 5902 4928
rect 5966 4864 5982 4928
rect 6046 4864 6062 4928
rect 6126 4864 6132 4928
rect 5816 4863 6132 4864
rect 7764 4928 8080 4929
rect 7764 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7930 4928
rect 7994 4864 8010 4928
rect 8074 4864 8080 4928
rect 7764 4863 8080 4864
rect 2894 4384 3210 4385
rect 2894 4320 2900 4384
rect 2964 4320 2980 4384
rect 3044 4320 3060 4384
rect 3124 4320 3140 4384
rect 3204 4320 3210 4384
rect 2894 4319 3210 4320
rect 4842 4384 5158 4385
rect 4842 4320 4848 4384
rect 4912 4320 4928 4384
rect 4992 4320 5008 4384
rect 5072 4320 5088 4384
rect 5152 4320 5158 4384
rect 4842 4319 5158 4320
rect 6790 4384 7106 4385
rect 6790 4320 6796 4384
rect 6860 4320 6876 4384
rect 6940 4320 6956 4384
rect 7020 4320 7036 4384
rect 7100 4320 7106 4384
rect 6790 4319 7106 4320
rect 1920 3840 2236 3841
rect 1920 3776 1926 3840
rect 1990 3776 2006 3840
rect 2070 3776 2086 3840
rect 2150 3776 2166 3840
rect 2230 3776 2236 3840
rect 1920 3775 2236 3776
rect 3868 3840 4184 3841
rect 3868 3776 3874 3840
rect 3938 3776 3954 3840
rect 4018 3776 4034 3840
rect 4098 3776 4114 3840
rect 4178 3776 4184 3840
rect 3868 3775 4184 3776
rect 5816 3840 6132 3841
rect 5816 3776 5822 3840
rect 5886 3776 5902 3840
rect 5966 3776 5982 3840
rect 6046 3776 6062 3840
rect 6126 3776 6132 3840
rect 5816 3775 6132 3776
rect 7764 3840 8080 3841
rect 7764 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7930 3840
rect 7994 3776 8010 3840
rect 8074 3776 8080 3840
rect 7764 3775 8080 3776
rect 2894 3296 3210 3297
rect 2894 3232 2900 3296
rect 2964 3232 2980 3296
rect 3044 3232 3060 3296
rect 3124 3232 3140 3296
rect 3204 3232 3210 3296
rect 2894 3231 3210 3232
rect 4842 3296 5158 3297
rect 4842 3232 4848 3296
rect 4912 3232 4928 3296
rect 4992 3232 5008 3296
rect 5072 3232 5088 3296
rect 5152 3232 5158 3296
rect 4842 3231 5158 3232
rect 6790 3296 7106 3297
rect 6790 3232 6796 3296
rect 6860 3232 6876 3296
rect 6940 3232 6956 3296
rect 7020 3232 7036 3296
rect 7100 3232 7106 3296
rect 6790 3231 7106 3232
rect 1920 2752 2236 2753
rect 1920 2688 1926 2752
rect 1990 2688 2006 2752
rect 2070 2688 2086 2752
rect 2150 2688 2166 2752
rect 2230 2688 2236 2752
rect 1920 2687 2236 2688
rect 3868 2752 4184 2753
rect 3868 2688 3874 2752
rect 3938 2688 3954 2752
rect 4018 2688 4034 2752
rect 4098 2688 4114 2752
rect 4178 2688 4184 2752
rect 3868 2687 4184 2688
rect 5816 2752 6132 2753
rect 5816 2688 5822 2752
rect 5886 2688 5902 2752
rect 5966 2688 5982 2752
rect 6046 2688 6062 2752
rect 6126 2688 6132 2752
rect 5816 2687 6132 2688
rect 7764 2752 8080 2753
rect 7764 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7930 2752
rect 7994 2688 8010 2752
rect 8074 2688 8080 2752
rect 7764 2687 8080 2688
rect 2894 2208 3210 2209
rect 2894 2144 2900 2208
rect 2964 2144 2980 2208
rect 3044 2144 3060 2208
rect 3124 2144 3140 2208
rect 3204 2144 3210 2208
rect 2894 2143 3210 2144
rect 4842 2208 5158 2209
rect 4842 2144 4848 2208
rect 4912 2144 4928 2208
rect 4992 2144 5008 2208
rect 5072 2144 5088 2208
rect 5152 2144 5158 2208
rect 4842 2143 5158 2144
rect 6790 2208 7106 2209
rect 6790 2144 6796 2208
rect 6860 2144 6876 2208
rect 6940 2144 6956 2208
rect 7020 2144 7036 2208
rect 7100 2144 7106 2208
rect 6790 2143 7106 2144
<< via3 >>
rect 2900 7644 2964 7648
rect 2900 7588 2904 7644
rect 2904 7588 2960 7644
rect 2960 7588 2964 7644
rect 2900 7584 2964 7588
rect 2980 7644 3044 7648
rect 2980 7588 2984 7644
rect 2984 7588 3040 7644
rect 3040 7588 3044 7644
rect 2980 7584 3044 7588
rect 3060 7644 3124 7648
rect 3060 7588 3064 7644
rect 3064 7588 3120 7644
rect 3120 7588 3124 7644
rect 3060 7584 3124 7588
rect 3140 7644 3204 7648
rect 3140 7588 3144 7644
rect 3144 7588 3200 7644
rect 3200 7588 3204 7644
rect 3140 7584 3204 7588
rect 4848 7644 4912 7648
rect 4848 7588 4852 7644
rect 4852 7588 4908 7644
rect 4908 7588 4912 7644
rect 4848 7584 4912 7588
rect 4928 7644 4992 7648
rect 4928 7588 4932 7644
rect 4932 7588 4988 7644
rect 4988 7588 4992 7644
rect 4928 7584 4992 7588
rect 5008 7644 5072 7648
rect 5008 7588 5012 7644
rect 5012 7588 5068 7644
rect 5068 7588 5072 7644
rect 5008 7584 5072 7588
rect 5088 7644 5152 7648
rect 5088 7588 5092 7644
rect 5092 7588 5148 7644
rect 5148 7588 5152 7644
rect 5088 7584 5152 7588
rect 6796 7644 6860 7648
rect 6796 7588 6800 7644
rect 6800 7588 6856 7644
rect 6856 7588 6860 7644
rect 6796 7584 6860 7588
rect 6876 7644 6940 7648
rect 6876 7588 6880 7644
rect 6880 7588 6936 7644
rect 6936 7588 6940 7644
rect 6876 7584 6940 7588
rect 6956 7644 7020 7648
rect 6956 7588 6960 7644
rect 6960 7588 7016 7644
rect 7016 7588 7020 7644
rect 6956 7584 7020 7588
rect 7036 7644 7100 7648
rect 7036 7588 7040 7644
rect 7040 7588 7096 7644
rect 7096 7588 7100 7644
rect 7036 7584 7100 7588
rect 1926 7100 1990 7104
rect 1926 7044 1930 7100
rect 1930 7044 1986 7100
rect 1986 7044 1990 7100
rect 1926 7040 1990 7044
rect 2006 7100 2070 7104
rect 2006 7044 2010 7100
rect 2010 7044 2066 7100
rect 2066 7044 2070 7100
rect 2006 7040 2070 7044
rect 2086 7100 2150 7104
rect 2086 7044 2090 7100
rect 2090 7044 2146 7100
rect 2146 7044 2150 7100
rect 2086 7040 2150 7044
rect 2166 7100 2230 7104
rect 2166 7044 2170 7100
rect 2170 7044 2226 7100
rect 2226 7044 2230 7100
rect 2166 7040 2230 7044
rect 3874 7100 3938 7104
rect 3874 7044 3878 7100
rect 3878 7044 3934 7100
rect 3934 7044 3938 7100
rect 3874 7040 3938 7044
rect 3954 7100 4018 7104
rect 3954 7044 3958 7100
rect 3958 7044 4014 7100
rect 4014 7044 4018 7100
rect 3954 7040 4018 7044
rect 4034 7100 4098 7104
rect 4034 7044 4038 7100
rect 4038 7044 4094 7100
rect 4094 7044 4098 7100
rect 4034 7040 4098 7044
rect 4114 7100 4178 7104
rect 4114 7044 4118 7100
rect 4118 7044 4174 7100
rect 4174 7044 4178 7100
rect 4114 7040 4178 7044
rect 5822 7100 5886 7104
rect 5822 7044 5826 7100
rect 5826 7044 5882 7100
rect 5882 7044 5886 7100
rect 5822 7040 5886 7044
rect 5902 7100 5966 7104
rect 5902 7044 5906 7100
rect 5906 7044 5962 7100
rect 5962 7044 5966 7100
rect 5902 7040 5966 7044
rect 5982 7100 6046 7104
rect 5982 7044 5986 7100
rect 5986 7044 6042 7100
rect 6042 7044 6046 7100
rect 5982 7040 6046 7044
rect 6062 7100 6126 7104
rect 6062 7044 6066 7100
rect 6066 7044 6122 7100
rect 6122 7044 6126 7100
rect 6062 7040 6126 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 7930 7100 7994 7104
rect 7930 7044 7934 7100
rect 7934 7044 7990 7100
rect 7990 7044 7994 7100
rect 7930 7040 7994 7044
rect 8010 7100 8074 7104
rect 8010 7044 8014 7100
rect 8014 7044 8070 7100
rect 8070 7044 8074 7100
rect 8010 7040 8074 7044
rect 2900 6556 2964 6560
rect 2900 6500 2904 6556
rect 2904 6500 2960 6556
rect 2960 6500 2964 6556
rect 2900 6496 2964 6500
rect 2980 6556 3044 6560
rect 2980 6500 2984 6556
rect 2984 6500 3040 6556
rect 3040 6500 3044 6556
rect 2980 6496 3044 6500
rect 3060 6556 3124 6560
rect 3060 6500 3064 6556
rect 3064 6500 3120 6556
rect 3120 6500 3124 6556
rect 3060 6496 3124 6500
rect 3140 6556 3204 6560
rect 3140 6500 3144 6556
rect 3144 6500 3200 6556
rect 3200 6500 3204 6556
rect 3140 6496 3204 6500
rect 4848 6556 4912 6560
rect 4848 6500 4852 6556
rect 4852 6500 4908 6556
rect 4908 6500 4912 6556
rect 4848 6496 4912 6500
rect 4928 6556 4992 6560
rect 4928 6500 4932 6556
rect 4932 6500 4988 6556
rect 4988 6500 4992 6556
rect 4928 6496 4992 6500
rect 5008 6556 5072 6560
rect 5008 6500 5012 6556
rect 5012 6500 5068 6556
rect 5068 6500 5072 6556
rect 5008 6496 5072 6500
rect 5088 6556 5152 6560
rect 5088 6500 5092 6556
rect 5092 6500 5148 6556
rect 5148 6500 5152 6556
rect 5088 6496 5152 6500
rect 6796 6556 6860 6560
rect 6796 6500 6800 6556
rect 6800 6500 6856 6556
rect 6856 6500 6860 6556
rect 6796 6496 6860 6500
rect 6876 6556 6940 6560
rect 6876 6500 6880 6556
rect 6880 6500 6936 6556
rect 6936 6500 6940 6556
rect 6876 6496 6940 6500
rect 6956 6556 7020 6560
rect 6956 6500 6960 6556
rect 6960 6500 7016 6556
rect 7016 6500 7020 6556
rect 6956 6496 7020 6500
rect 7036 6556 7100 6560
rect 7036 6500 7040 6556
rect 7040 6500 7096 6556
rect 7096 6500 7100 6556
rect 7036 6496 7100 6500
rect 1926 6012 1990 6016
rect 1926 5956 1930 6012
rect 1930 5956 1986 6012
rect 1986 5956 1990 6012
rect 1926 5952 1990 5956
rect 2006 6012 2070 6016
rect 2006 5956 2010 6012
rect 2010 5956 2066 6012
rect 2066 5956 2070 6012
rect 2006 5952 2070 5956
rect 2086 6012 2150 6016
rect 2086 5956 2090 6012
rect 2090 5956 2146 6012
rect 2146 5956 2150 6012
rect 2086 5952 2150 5956
rect 2166 6012 2230 6016
rect 2166 5956 2170 6012
rect 2170 5956 2226 6012
rect 2226 5956 2230 6012
rect 2166 5952 2230 5956
rect 3874 6012 3938 6016
rect 3874 5956 3878 6012
rect 3878 5956 3934 6012
rect 3934 5956 3938 6012
rect 3874 5952 3938 5956
rect 3954 6012 4018 6016
rect 3954 5956 3958 6012
rect 3958 5956 4014 6012
rect 4014 5956 4018 6012
rect 3954 5952 4018 5956
rect 4034 6012 4098 6016
rect 4034 5956 4038 6012
rect 4038 5956 4094 6012
rect 4094 5956 4098 6012
rect 4034 5952 4098 5956
rect 4114 6012 4178 6016
rect 4114 5956 4118 6012
rect 4118 5956 4174 6012
rect 4174 5956 4178 6012
rect 4114 5952 4178 5956
rect 5822 6012 5886 6016
rect 5822 5956 5826 6012
rect 5826 5956 5882 6012
rect 5882 5956 5886 6012
rect 5822 5952 5886 5956
rect 5902 6012 5966 6016
rect 5902 5956 5906 6012
rect 5906 5956 5962 6012
rect 5962 5956 5966 6012
rect 5902 5952 5966 5956
rect 5982 6012 6046 6016
rect 5982 5956 5986 6012
rect 5986 5956 6042 6012
rect 6042 5956 6046 6012
rect 5982 5952 6046 5956
rect 6062 6012 6126 6016
rect 6062 5956 6066 6012
rect 6066 5956 6122 6012
rect 6122 5956 6126 6012
rect 6062 5952 6126 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 7930 6012 7994 6016
rect 7930 5956 7934 6012
rect 7934 5956 7990 6012
rect 7990 5956 7994 6012
rect 7930 5952 7994 5956
rect 8010 6012 8074 6016
rect 8010 5956 8014 6012
rect 8014 5956 8070 6012
rect 8070 5956 8074 6012
rect 8010 5952 8074 5956
rect 2900 5468 2964 5472
rect 2900 5412 2904 5468
rect 2904 5412 2960 5468
rect 2960 5412 2964 5468
rect 2900 5408 2964 5412
rect 2980 5468 3044 5472
rect 2980 5412 2984 5468
rect 2984 5412 3040 5468
rect 3040 5412 3044 5468
rect 2980 5408 3044 5412
rect 3060 5468 3124 5472
rect 3060 5412 3064 5468
rect 3064 5412 3120 5468
rect 3120 5412 3124 5468
rect 3060 5408 3124 5412
rect 3140 5468 3204 5472
rect 3140 5412 3144 5468
rect 3144 5412 3200 5468
rect 3200 5412 3204 5468
rect 3140 5408 3204 5412
rect 4848 5468 4912 5472
rect 4848 5412 4852 5468
rect 4852 5412 4908 5468
rect 4908 5412 4912 5468
rect 4848 5408 4912 5412
rect 4928 5468 4992 5472
rect 4928 5412 4932 5468
rect 4932 5412 4988 5468
rect 4988 5412 4992 5468
rect 4928 5408 4992 5412
rect 5008 5468 5072 5472
rect 5008 5412 5012 5468
rect 5012 5412 5068 5468
rect 5068 5412 5072 5468
rect 5008 5408 5072 5412
rect 5088 5468 5152 5472
rect 5088 5412 5092 5468
rect 5092 5412 5148 5468
rect 5148 5412 5152 5468
rect 5088 5408 5152 5412
rect 6796 5468 6860 5472
rect 6796 5412 6800 5468
rect 6800 5412 6856 5468
rect 6856 5412 6860 5468
rect 6796 5408 6860 5412
rect 6876 5468 6940 5472
rect 6876 5412 6880 5468
rect 6880 5412 6936 5468
rect 6936 5412 6940 5468
rect 6876 5408 6940 5412
rect 6956 5468 7020 5472
rect 6956 5412 6960 5468
rect 6960 5412 7016 5468
rect 7016 5412 7020 5468
rect 6956 5408 7020 5412
rect 7036 5468 7100 5472
rect 7036 5412 7040 5468
rect 7040 5412 7096 5468
rect 7096 5412 7100 5468
rect 7036 5408 7100 5412
rect 1926 4924 1990 4928
rect 1926 4868 1930 4924
rect 1930 4868 1986 4924
rect 1986 4868 1990 4924
rect 1926 4864 1990 4868
rect 2006 4924 2070 4928
rect 2006 4868 2010 4924
rect 2010 4868 2066 4924
rect 2066 4868 2070 4924
rect 2006 4864 2070 4868
rect 2086 4924 2150 4928
rect 2086 4868 2090 4924
rect 2090 4868 2146 4924
rect 2146 4868 2150 4924
rect 2086 4864 2150 4868
rect 2166 4924 2230 4928
rect 2166 4868 2170 4924
rect 2170 4868 2226 4924
rect 2226 4868 2230 4924
rect 2166 4864 2230 4868
rect 3874 4924 3938 4928
rect 3874 4868 3878 4924
rect 3878 4868 3934 4924
rect 3934 4868 3938 4924
rect 3874 4864 3938 4868
rect 3954 4924 4018 4928
rect 3954 4868 3958 4924
rect 3958 4868 4014 4924
rect 4014 4868 4018 4924
rect 3954 4864 4018 4868
rect 4034 4924 4098 4928
rect 4034 4868 4038 4924
rect 4038 4868 4094 4924
rect 4094 4868 4098 4924
rect 4034 4864 4098 4868
rect 4114 4924 4178 4928
rect 4114 4868 4118 4924
rect 4118 4868 4174 4924
rect 4174 4868 4178 4924
rect 4114 4864 4178 4868
rect 5822 4924 5886 4928
rect 5822 4868 5826 4924
rect 5826 4868 5882 4924
rect 5882 4868 5886 4924
rect 5822 4864 5886 4868
rect 5902 4924 5966 4928
rect 5902 4868 5906 4924
rect 5906 4868 5962 4924
rect 5962 4868 5966 4924
rect 5902 4864 5966 4868
rect 5982 4924 6046 4928
rect 5982 4868 5986 4924
rect 5986 4868 6042 4924
rect 6042 4868 6046 4924
rect 5982 4864 6046 4868
rect 6062 4924 6126 4928
rect 6062 4868 6066 4924
rect 6066 4868 6122 4924
rect 6122 4868 6126 4924
rect 6062 4864 6126 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 7930 4924 7994 4928
rect 7930 4868 7934 4924
rect 7934 4868 7990 4924
rect 7990 4868 7994 4924
rect 7930 4864 7994 4868
rect 8010 4924 8074 4928
rect 8010 4868 8014 4924
rect 8014 4868 8070 4924
rect 8070 4868 8074 4924
rect 8010 4864 8074 4868
rect 2900 4380 2964 4384
rect 2900 4324 2904 4380
rect 2904 4324 2960 4380
rect 2960 4324 2964 4380
rect 2900 4320 2964 4324
rect 2980 4380 3044 4384
rect 2980 4324 2984 4380
rect 2984 4324 3040 4380
rect 3040 4324 3044 4380
rect 2980 4320 3044 4324
rect 3060 4380 3124 4384
rect 3060 4324 3064 4380
rect 3064 4324 3120 4380
rect 3120 4324 3124 4380
rect 3060 4320 3124 4324
rect 3140 4380 3204 4384
rect 3140 4324 3144 4380
rect 3144 4324 3200 4380
rect 3200 4324 3204 4380
rect 3140 4320 3204 4324
rect 4848 4380 4912 4384
rect 4848 4324 4852 4380
rect 4852 4324 4908 4380
rect 4908 4324 4912 4380
rect 4848 4320 4912 4324
rect 4928 4380 4992 4384
rect 4928 4324 4932 4380
rect 4932 4324 4988 4380
rect 4988 4324 4992 4380
rect 4928 4320 4992 4324
rect 5008 4380 5072 4384
rect 5008 4324 5012 4380
rect 5012 4324 5068 4380
rect 5068 4324 5072 4380
rect 5008 4320 5072 4324
rect 5088 4380 5152 4384
rect 5088 4324 5092 4380
rect 5092 4324 5148 4380
rect 5148 4324 5152 4380
rect 5088 4320 5152 4324
rect 6796 4380 6860 4384
rect 6796 4324 6800 4380
rect 6800 4324 6856 4380
rect 6856 4324 6860 4380
rect 6796 4320 6860 4324
rect 6876 4380 6940 4384
rect 6876 4324 6880 4380
rect 6880 4324 6936 4380
rect 6936 4324 6940 4380
rect 6876 4320 6940 4324
rect 6956 4380 7020 4384
rect 6956 4324 6960 4380
rect 6960 4324 7016 4380
rect 7016 4324 7020 4380
rect 6956 4320 7020 4324
rect 7036 4380 7100 4384
rect 7036 4324 7040 4380
rect 7040 4324 7096 4380
rect 7096 4324 7100 4380
rect 7036 4320 7100 4324
rect 1926 3836 1990 3840
rect 1926 3780 1930 3836
rect 1930 3780 1986 3836
rect 1986 3780 1990 3836
rect 1926 3776 1990 3780
rect 2006 3836 2070 3840
rect 2006 3780 2010 3836
rect 2010 3780 2066 3836
rect 2066 3780 2070 3836
rect 2006 3776 2070 3780
rect 2086 3836 2150 3840
rect 2086 3780 2090 3836
rect 2090 3780 2146 3836
rect 2146 3780 2150 3836
rect 2086 3776 2150 3780
rect 2166 3836 2230 3840
rect 2166 3780 2170 3836
rect 2170 3780 2226 3836
rect 2226 3780 2230 3836
rect 2166 3776 2230 3780
rect 3874 3836 3938 3840
rect 3874 3780 3878 3836
rect 3878 3780 3934 3836
rect 3934 3780 3938 3836
rect 3874 3776 3938 3780
rect 3954 3836 4018 3840
rect 3954 3780 3958 3836
rect 3958 3780 4014 3836
rect 4014 3780 4018 3836
rect 3954 3776 4018 3780
rect 4034 3836 4098 3840
rect 4034 3780 4038 3836
rect 4038 3780 4094 3836
rect 4094 3780 4098 3836
rect 4034 3776 4098 3780
rect 4114 3836 4178 3840
rect 4114 3780 4118 3836
rect 4118 3780 4174 3836
rect 4174 3780 4178 3836
rect 4114 3776 4178 3780
rect 5822 3836 5886 3840
rect 5822 3780 5826 3836
rect 5826 3780 5882 3836
rect 5882 3780 5886 3836
rect 5822 3776 5886 3780
rect 5902 3836 5966 3840
rect 5902 3780 5906 3836
rect 5906 3780 5962 3836
rect 5962 3780 5966 3836
rect 5902 3776 5966 3780
rect 5982 3836 6046 3840
rect 5982 3780 5986 3836
rect 5986 3780 6042 3836
rect 6042 3780 6046 3836
rect 5982 3776 6046 3780
rect 6062 3836 6126 3840
rect 6062 3780 6066 3836
rect 6066 3780 6122 3836
rect 6122 3780 6126 3836
rect 6062 3776 6126 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 7930 3836 7994 3840
rect 7930 3780 7934 3836
rect 7934 3780 7990 3836
rect 7990 3780 7994 3836
rect 7930 3776 7994 3780
rect 8010 3836 8074 3840
rect 8010 3780 8014 3836
rect 8014 3780 8070 3836
rect 8070 3780 8074 3836
rect 8010 3776 8074 3780
rect 2900 3292 2964 3296
rect 2900 3236 2904 3292
rect 2904 3236 2960 3292
rect 2960 3236 2964 3292
rect 2900 3232 2964 3236
rect 2980 3292 3044 3296
rect 2980 3236 2984 3292
rect 2984 3236 3040 3292
rect 3040 3236 3044 3292
rect 2980 3232 3044 3236
rect 3060 3292 3124 3296
rect 3060 3236 3064 3292
rect 3064 3236 3120 3292
rect 3120 3236 3124 3292
rect 3060 3232 3124 3236
rect 3140 3292 3204 3296
rect 3140 3236 3144 3292
rect 3144 3236 3200 3292
rect 3200 3236 3204 3292
rect 3140 3232 3204 3236
rect 4848 3292 4912 3296
rect 4848 3236 4852 3292
rect 4852 3236 4908 3292
rect 4908 3236 4912 3292
rect 4848 3232 4912 3236
rect 4928 3292 4992 3296
rect 4928 3236 4932 3292
rect 4932 3236 4988 3292
rect 4988 3236 4992 3292
rect 4928 3232 4992 3236
rect 5008 3292 5072 3296
rect 5008 3236 5012 3292
rect 5012 3236 5068 3292
rect 5068 3236 5072 3292
rect 5008 3232 5072 3236
rect 5088 3292 5152 3296
rect 5088 3236 5092 3292
rect 5092 3236 5148 3292
rect 5148 3236 5152 3292
rect 5088 3232 5152 3236
rect 6796 3292 6860 3296
rect 6796 3236 6800 3292
rect 6800 3236 6856 3292
rect 6856 3236 6860 3292
rect 6796 3232 6860 3236
rect 6876 3292 6940 3296
rect 6876 3236 6880 3292
rect 6880 3236 6936 3292
rect 6936 3236 6940 3292
rect 6876 3232 6940 3236
rect 6956 3292 7020 3296
rect 6956 3236 6960 3292
rect 6960 3236 7016 3292
rect 7016 3236 7020 3292
rect 6956 3232 7020 3236
rect 7036 3292 7100 3296
rect 7036 3236 7040 3292
rect 7040 3236 7096 3292
rect 7096 3236 7100 3292
rect 7036 3232 7100 3236
rect 1926 2748 1990 2752
rect 1926 2692 1930 2748
rect 1930 2692 1986 2748
rect 1986 2692 1990 2748
rect 1926 2688 1990 2692
rect 2006 2748 2070 2752
rect 2006 2692 2010 2748
rect 2010 2692 2066 2748
rect 2066 2692 2070 2748
rect 2006 2688 2070 2692
rect 2086 2748 2150 2752
rect 2086 2692 2090 2748
rect 2090 2692 2146 2748
rect 2146 2692 2150 2748
rect 2086 2688 2150 2692
rect 2166 2748 2230 2752
rect 2166 2692 2170 2748
rect 2170 2692 2226 2748
rect 2226 2692 2230 2748
rect 2166 2688 2230 2692
rect 3874 2748 3938 2752
rect 3874 2692 3878 2748
rect 3878 2692 3934 2748
rect 3934 2692 3938 2748
rect 3874 2688 3938 2692
rect 3954 2748 4018 2752
rect 3954 2692 3958 2748
rect 3958 2692 4014 2748
rect 4014 2692 4018 2748
rect 3954 2688 4018 2692
rect 4034 2748 4098 2752
rect 4034 2692 4038 2748
rect 4038 2692 4094 2748
rect 4094 2692 4098 2748
rect 4034 2688 4098 2692
rect 4114 2748 4178 2752
rect 4114 2692 4118 2748
rect 4118 2692 4174 2748
rect 4174 2692 4178 2748
rect 4114 2688 4178 2692
rect 5822 2748 5886 2752
rect 5822 2692 5826 2748
rect 5826 2692 5882 2748
rect 5882 2692 5886 2748
rect 5822 2688 5886 2692
rect 5902 2748 5966 2752
rect 5902 2692 5906 2748
rect 5906 2692 5962 2748
rect 5962 2692 5966 2748
rect 5902 2688 5966 2692
rect 5982 2748 6046 2752
rect 5982 2692 5986 2748
rect 5986 2692 6042 2748
rect 6042 2692 6046 2748
rect 5982 2688 6046 2692
rect 6062 2748 6126 2752
rect 6062 2692 6066 2748
rect 6066 2692 6122 2748
rect 6122 2692 6126 2748
rect 6062 2688 6126 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 7930 2748 7994 2752
rect 7930 2692 7934 2748
rect 7934 2692 7990 2748
rect 7990 2692 7994 2748
rect 7930 2688 7994 2692
rect 8010 2748 8074 2752
rect 8010 2692 8014 2748
rect 8014 2692 8070 2748
rect 8070 2692 8074 2748
rect 8010 2688 8074 2692
rect 2900 2204 2964 2208
rect 2900 2148 2904 2204
rect 2904 2148 2960 2204
rect 2960 2148 2964 2204
rect 2900 2144 2964 2148
rect 2980 2204 3044 2208
rect 2980 2148 2984 2204
rect 2984 2148 3040 2204
rect 3040 2148 3044 2204
rect 2980 2144 3044 2148
rect 3060 2204 3124 2208
rect 3060 2148 3064 2204
rect 3064 2148 3120 2204
rect 3120 2148 3124 2204
rect 3060 2144 3124 2148
rect 3140 2204 3204 2208
rect 3140 2148 3144 2204
rect 3144 2148 3200 2204
rect 3200 2148 3204 2204
rect 3140 2144 3204 2148
rect 4848 2204 4912 2208
rect 4848 2148 4852 2204
rect 4852 2148 4908 2204
rect 4908 2148 4912 2204
rect 4848 2144 4912 2148
rect 4928 2204 4992 2208
rect 4928 2148 4932 2204
rect 4932 2148 4988 2204
rect 4988 2148 4992 2204
rect 4928 2144 4992 2148
rect 5008 2204 5072 2208
rect 5008 2148 5012 2204
rect 5012 2148 5068 2204
rect 5068 2148 5072 2204
rect 5008 2144 5072 2148
rect 5088 2204 5152 2208
rect 5088 2148 5092 2204
rect 5092 2148 5148 2204
rect 5148 2148 5152 2204
rect 5088 2144 5152 2148
rect 6796 2204 6860 2208
rect 6796 2148 6800 2204
rect 6800 2148 6856 2204
rect 6856 2148 6860 2204
rect 6796 2144 6860 2148
rect 6876 2204 6940 2208
rect 6876 2148 6880 2204
rect 6880 2148 6936 2204
rect 6936 2148 6940 2204
rect 6876 2144 6940 2148
rect 6956 2204 7020 2208
rect 6956 2148 6960 2204
rect 6960 2148 7016 2204
rect 7016 2148 7020 2204
rect 6956 2144 7020 2148
rect 7036 2204 7100 2208
rect 7036 2148 7040 2204
rect 7040 2148 7096 2204
rect 7096 2148 7100 2204
rect 7036 2144 7100 2148
<< metal4 >>
rect 1918 7104 2238 7664
rect 1918 7040 1926 7104
rect 1990 7040 2006 7104
rect 2070 7040 2086 7104
rect 2150 7040 2166 7104
rect 2230 7040 2238 7104
rect 1918 6016 2238 7040
rect 1918 5952 1926 6016
rect 1990 5952 2006 6016
rect 2070 5952 2086 6016
rect 2150 5952 2166 6016
rect 2230 5952 2238 6016
rect 1918 4928 2238 5952
rect 1918 4864 1926 4928
rect 1990 4864 2006 4928
rect 2070 4864 2086 4928
rect 2150 4864 2166 4928
rect 2230 4864 2238 4928
rect 1918 3840 2238 4864
rect 1918 3776 1926 3840
rect 1990 3776 2006 3840
rect 2070 3776 2086 3840
rect 2150 3776 2166 3840
rect 2230 3776 2238 3840
rect 1918 2752 2238 3776
rect 1918 2688 1926 2752
rect 1990 2688 2006 2752
rect 2070 2688 2086 2752
rect 2150 2688 2166 2752
rect 2230 2688 2238 2752
rect 1918 2128 2238 2688
rect 2892 7648 3212 7664
rect 2892 7584 2900 7648
rect 2964 7584 2980 7648
rect 3044 7584 3060 7648
rect 3124 7584 3140 7648
rect 3204 7584 3212 7648
rect 2892 6560 3212 7584
rect 2892 6496 2900 6560
rect 2964 6496 2980 6560
rect 3044 6496 3060 6560
rect 3124 6496 3140 6560
rect 3204 6496 3212 6560
rect 2892 5472 3212 6496
rect 2892 5408 2900 5472
rect 2964 5408 2980 5472
rect 3044 5408 3060 5472
rect 3124 5408 3140 5472
rect 3204 5408 3212 5472
rect 2892 4384 3212 5408
rect 2892 4320 2900 4384
rect 2964 4320 2980 4384
rect 3044 4320 3060 4384
rect 3124 4320 3140 4384
rect 3204 4320 3212 4384
rect 2892 3296 3212 4320
rect 2892 3232 2900 3296
rect 2964 3232 2980 3296
rect 3044 3232 3060 3296
rect 3124 3232 3140 3296
rect 3204 3232 3212 3296
rect 2892 2208 3212 3232
rect 2892 2144 2900 2208
rect 2964 2144 2980 2208
rect 3044 2144 3060 2208
rect 3124 2144 3140 2208
rect 3204 2144 3212 2208
rect 2892 2128 3212 2144
rect 3866 7104 4186 7664
rect 3866 7040 3874 7104
rect 3938 7040 3954 7104
rect 4018 7040 4034 7104
rect 4098 7040 4114 7104
rect 4178 7040 4186 7104
rect 3866 6016 4186 7040
rect 3866 5952 3874 6016
rect 3938 5952 3954 6016
rect 4018 5952 4034 6016
rect 4098 5952 4114 6016
rect 4178 5952 4186 6016
rect 3866 4928 4186 5952
rect 3866 4864 3874 4928
rect 3938 4864 3954 4928
rect 4018 4864 4034 4928
rect 4098 4864 4114 4928
rect 4178 4864 4186 4928
rect 3866 3840 4186 4864
rect 3866 3776 3874 3840
rect 3938 3776 3954 3840
rect 4018 3776 4034 3840
rect 4098 3776 4114 3840
rect 4178 3776 4186 3840
rect 3866 2752 4186 3776
rect 3866 2688 3874 2752
rect 3938 2688 3954 2752
rect 4018 2688 4034 2752
rect 4098 2688 4114 2752
rect 4178 2688 4186 2752
rect 3866 2128 4186 2688
rect 4840 7648 5160 7664
rect 4840 7584 4848 7648
rect 4912 7584 4928 7648
rect 4992 7584 5008 7648
rect 5072 7584 5088 7648
rect 5152 7584 5160 7648
rect 4840 6560 5160 7584
rect 4840 6496 4848 6560
rect 4912 6496 4928 6560
rect 4992 6496 5008 6560
rect 5072 6496 5088 6560
rect 5152 6496 5160 6560
rect 4840 5472 5160 6496
rect 4840 5408 4848 5472
rect 4912 5408 4928 5472
rect 4992 5408 5008 5472
rect 5072 5408 5088 5472
rect 5152 5408 5160 5472
rect 4840 4384 5160 5408
rect 4840 4320 4848 4384
rect 4912 4320 4928 4384
rect 4992 4320 5008 4384
rect 5072 4320 5088 4384
rect 5152 4320 5160 4384
rect 4840 3296 5160 4320
rect 4840 3232 4848 3296
rect 4912 3232 4928 3296
rect 4992 3232 5008 3296
rect 5072 3232 5088 3296
rect 5152 3232 5160 3296
rect 4840 2208 5160 3232
rect 4840 2144 4848 2208
rect 4912 2144 4928 2208
rect 4992 2144 5008 2208
rect 5072 2144 5088 2208
rect 5152 2144 5160 2208
rect 4840 2128 5160 2144
rect 5814 7104 6134 7664
rect 5814 7040 5822 7104
rect 5886 7040 5902 7104
rect 5966 7040 5982 7104
rect 6046 7040 6062 7104
rect 6126 7040 6134 7104
rect 5814 6016 6134 7040
rect 5814 5952 5822 6016
rect 5886 5952 5902 6016
rect 5966 5952 5982 6016
rect 6046 5952 6062 6016
rect 6126 5952 6134 6016
rect 5814 4928 6134 5952
rect 5814 4864 5822 4928
rect 5886 4864 5902 4928
rect 5966 4864 5982 4928
rect 6046 4864 6062 4928
rect 6126 4864 6134 4928
rect 5814 3840 6134 4864
rect 5814 3776 5822 3840
rect 5886 3776 5902 3840
rect 5966 3776 5982 3840
rect 6046 3776 6062 3840
rect 6126 3776 6134 3840
rect 5814 2752 6134 3776
rect 5814 2688 5822 2752
rect 5886 2688 5902 2752
rect 5966 2688 5982 2752
rect 6046 2688 6062 2752
rect 6126 2688 6134 2752
rect 5814 2128 6134 2688
rect 6788 7648 7108 7664
rect 6788 7584 6796 7648
rect 6860 7584 6876 7648
rect 6940 7584 6956 7648
rect 7020 7584 7036 7648
rect 7100 7584 7108 7648
rect 6788 6560 7108 7584
rect 6788 6496 6796 6560
rect 6860 6496 6876 6560
rect 6940 6496 6956 6560
rect 7020 6496 7036 6560
rect 7100 6496 7108 6560
rect 6788 5472 7108 6496
rect 6788 5408 6796 5472
rect 6860 5408 6876 5472
rect 6940 5408 6956 5472
rect 7020 5408 7036 5472
rect 7100 5408 7108 5472
rect 6788 4384 7108 5408
rect 6788 4320 6796 4384
rect 6860 4320 6876 4384
rect 6940 4320 6956 4384
rect 7020 4320 7036 4384
rect 7100 4320 7108 4384
rect 6788 3296 7108 4320
rect 6788 3232 6796 3296
rect 6860 3232 6876 3296
rect 6940 3232 6956 3296
rect 7020 3232 7036 3296
rect 7100 3232 7108 3296
rect 6788 2208 7108 3232
rect 6788 2144 6796 2208
rect 6860 2144 6876 2208
rect 6940 2144 6956 2208
rect 7020 2144 7036 2208
rect 7100 2144 7108 2208
rect 6788 2128 7108 2144
rect 7762 7104 8082 7664
rect 7762 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7930 7104
rect 7994 7040 8010 7104
rect 8074 7040 8082 7104
rect 7762 6016 8082 7040
rect 7762 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7930 6016
rect 7994 5952 8010 6016
rect 8074 5952 8082 6016
rect 7762 4928 8082 5952
rect 7762 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7930 4928
rect 7994 4864 8010 4928
rect 8074 4864 8082 4928
rect 7762 3840 8082 4864
rect 7762 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7930 3840
rect 7994 3776 8010 3840
rect 8074 3776 8082 3840
rect 7762 2752 8082 3776
rect 7762 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7930 2752
rect 7994 2688 8010 2752
rect 8074 2688 8082 2752
rect 7762 2128 8082 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 8188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_55
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_67
timestamp 1649977179
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1649977179
transform 1 0 8372 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_64
timestamp 1649977179
transform 1 0 6992 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1649977179
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1649977179
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1649977179
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_75
timestamp 1649977179
transform 1 0 8004 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_42
timestamp 1649977179
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1649977179
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_70
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_62
timestamp 1649977179
transform 1 0 6808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_74
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1649977179
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1649977179
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1649977179
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _10_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _11_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _12_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _13_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _14_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _15_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _16_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _17_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _18_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _19_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6992 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1649977179
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _21_
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _22_
timestamp 1649977179
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _23_
timestamp 1649977179
transform -1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _24_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4324 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _25_
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _26_
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8188 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
<< labels >>
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clock
port 0 nsew signal input
flabel metal2 s 18 9200 74 10000 0 FreeSans 224 90 0 0 detector_out
port 1 nsew signal tristate
flabel metal2 s 9678 9200 9734 10000 0 FreeSans 224 90 0 0 reset
port 2 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 sequence_in
port 3 nsew signal input
flabel metal4 s 1918 2128 2238 7664 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 3866 2128 4186 7664 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 5814 2128 6134 7664 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 7762 2128 8082 7664 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 2892 2128 3212 7664 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal4 s 4840 2128 5160 7664 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal4 s 6788 2128 7108 7664 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
